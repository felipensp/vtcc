@[translated]
module lib

@[export: 'tcc_backtrace']
pub fn tcc_backtrace(fmt &char) int {
	return 0
}
