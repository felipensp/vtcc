@[translated]
module lib

pub fn tcc_backtrace(fmt &char) {
}
