@[translated]
module main

@[hidden]
__global __dso_handle = unsafe { nil }
