@[translated]
module main

fn preprocess(is_bof int)  {
	s1 := tcc_state
	i := 0
	c := 0
	n := 0
	saved_parse_flags := 0
	
	buf := [1024]i8{}
	q := &i8(0)
	
	s := &Sym(0)
	saved_parse_flags = parse_flags
	parse_flags = 1 | 2 | 64 | 4 | (parse_flags & 8)
	next_nomacro()
	// RRRREG redo id=0x7fffc1b2a548
	redo: 
	match (tok) {
	 .tok_define{ // case comp body kind=BinaryOperator is_enum=true
	pp_debug_tok = tok
	next_nomacro()
	pp_debug_symv = tok
	parse_define()
	
	}
	 .tok_undef{ // case comp body kind=BinaryOperator is_enum=true
	pp_debug_tok = tok
	next_nomacro()
	pp_debug_symv = tok
	s = define_find(tok)
	if s {
	define_undef(s)
	}
	
	}
	 .tok_include, .tok_include_next{
	ch = file.buf_ptr [0] 
	skip_spaces()
	if ch == `<` {
		c = `>`
		goto read_name // id: 0x7fffc1b23c08
	}
	else if ch == `"` {
		c = ch
		// RRRREG read_name id=0x7fffc1b23c08
		read_name: 
		inp()
		q = buf
		for ch != c && ch != `\n` && ch != (-1) {
			if (q - buf) < sizeof(buf) - 1 {
			*q ++ = ch
			}
			if ch == `\\` {
				if handle_stray_noerror() == 0 {
				q --$
				}
			}
			else { // 3
			inp()
}
		}
		*q = ` `
		minp()
	}
	else {
		len := 0
		parse_flags = (1 | 4 | (parse_flags & 8))
		next()
		buf [0]  = ` `
		for tok != 10 {
			pstrcat(buf, sizeof(buf), get_tok_str(tok, &tokc))
			next()
		}
		len = C.strlen(buf)
		if (len < 2 || ((buf [0]  != `"` || buf [len - 1]  != `"`) && (buf [0]  != `<` || buf [len - 1]  != `>`))) {
		tcc_error(c"'#include' expects \"FILENAME\" or <FILENAME>")
		}
		c = buf [len - 1] 
		C.memmove(buf, buf + 1, len - 2)
		buf [len - 2]  = ` `
	}
	if s1.include_stack_ptr >= s1.include_stack + 32 {
	tcc_error(c'#include recursion too deep')
	}
	*s1.include_stack_ptr ++ = file
	i = if tok == Tcc_token.tok_include_next{ file.include_next_index } else {0}
	n = 2 + s1.nb_include_paths + s1.nb_sysinclude_paths
	for  ; i < n ; i ++ {
		buf1 := [1024]i8{}
		e := &CachedInclude(0)
		path := &i8(0)
		if i == 0 {
			if !(buf [0]  == `/`) {
			continue
			
			}
			buf1 [0]  = 0
		}
		else if i == 1 {
			if c != `"` {
			continue
			
			}
			path = file.truefilename
			pstrncpy(buf1, path, tcc_basename(path) - path)
		}
		else {
			j := i - 2
k := j - s1.nb_include_paths

			path = if k < 0{ s1.include_paths [j]  } else {s1.sysinclude_paths [k] }
			pstrcpy(buf1, sizeof(buf1), path)
			pstrcat(buf1, sizeof(buf1), c'/')
		}
		pstrcat(buf1, sizeof(buf1), buf)
		e = search_cached_include(s1, buf1, 0)
		if e && (define_find(e.ifndef_macro) || e.once == pp_once) {
			goto include_done // id: 0x7fffc1b27880
		}
		if tcc_open(s1, buf1) < 0 {
		continue
		
		}
		file.include_next_index = i + 1
		if s1.gen_deps {
			dynarray_add(&s1.target_deps, &s1.nb_target_deps, tcc_strdup(buf1))
		}
		if s1.do_debug {
		put_stabs(file.filename, __stab_debug_code.n_bincl, 0, 0, 0)
		}
		tok_flags |= 2 | 1
		ch = file.buf_ptr [0] 
		goto _GOTO_PLACEHOLDER_0x7fffc1b28330 // id: 0x7fffc1b28330
	}
	tcc_error(c"include file '%s' not found", buf)
	// RRRREG include_done id=0x7fffc1b27880
	include_done: 
	s1.include_stack_ptr --$
	
	}
	 .tok_ifndef{ // case comp body kind=BinaryOperator is_enum=true
	c = 1
	goto do_ifdef // id: 0x7fffc1b286c0
	}
	 .tok_if{ // case comp body kind=BinaryOperator is_enum=true
	c = expr_preprocess()
	goto do_if // id: 0x7fffc1b28820
	}
	 .tok_ifdef{ // case comp body kind=BinaryOperator is_enum=true
	c = 0
	// RRRREG do_ifdef id=0x7fffc1b286c0
	do_ifdef: 
	next_nomacro()
	if tok < 256 {
	tcc_error(c"invalid argument for '#if%sdef'", if c{ c'n' } else {c''})
	}
	if is_bof {
		if c {
			file.ifndef_macro = tok
		}
	}
	c = (define_find(tok) != 0) ^ c
	// RRRREG do_if id=0x7fffc1b28820
	do_if: 
	if s1.ifdef_stack_ptr >= s1.ifdef_stack + 64 {
	tcc_error(c'memory full (ifdef)')
	}
	*s1.ifdef_stack_ptr ++ = c
	goto test_skip // id: 0x7fffc1b29290
	}
	 .tok_else{ // case comp body kind=IfStmt is_enum=true
	if s1.ifdef_stack_ptr == s1.ifdef_stack {
	tcc_error(c'#else without matching #if')
	}
	if s1.ifdef_stack_ptr [-1]  & 2 {
	tcc_error(c'#else after #else')
	}
	c = (s1.ifdef_stack_ptr [-1]  ^= 3)
	goto test_else // id: 0x7fffc1b29938
	}
	 .tok_elif{ // case comp body kind=IfStmt is_enum=true
	if s1.ifdef_stack_ptr == s1.ifdef_stack {
	tcc_error(c'#elif without matching #if')
	}
	c = s1.ifdef_stack_ptr [-1] 
	if c > 1 {
	tcc_error(c'#elif after #else')
	}
	if c == 1 {
		c = 0
	}
	else {
		c = expr_preprocess()
		s1.ifdef_stack_ptr [-1]  = c
	}
	// RRRREG test_else id=0x7fffc1b29938
	test_else: 
	if s1.ifdef_stack_ptr == file.ifdef_stack_ptr + 1 {
	file.ifndef_macro = 0
	}
	// RRRREG test_skip id=0x7fffc1b29290
	test_skip: 
	if !(c & 1) {
		preprocess_skip()
		is_bof = 0
		goto _GOTO_PLACEHOLDER_0x7fffc1b2a548 // id: 0x7fffc1b2a548
	}
	
	}
	 .tok_endif{ // case comp body kind=IfStmt is_enum=true
	if s1.ifdef_stack_ptr <= file.ifdef_stack_ptr {
	tcc_error(c'#endif without matching #if')
	}
	s1.ifdef_stack_ptr --
	if file.ifndef_macro && s1.ifdef_stack_ptr == file.ifdef_stack_ptr {
		file.ifndef_macro_saved = file.ifndef_macro
		file.ifndef_macro = 0
		for tok != 10 {
		next_nomacro()
		}
		tok_flags |= 4
		goto _GOTO_PLACEHOLDER_0x7fffc1b28330 // id: 0x7fffc1b28330
	}
	
	}
	 190{ // case comp body kind=BinaryOperator is_enum=true
	n = strtoul(&i8(tokc.str.data), &q, 10)
	goto _line_num // id: 0x7fffc1b2b0e8
	}
	 .tok_line{ // case comp body kind=CallExpr is_enum=true
	next()
	if tok != 181 {
	// RRRREG _line_err id=0x7fffc1b2d3a8
	_line_err: 
	tcc_error(c'wrong #line format')
	}
	n = tokc.i
	// RRRREG _line_num id=0x7fffc1b2b0e8
	_line_num: 
	next()
	if tok != 10 {
		if tok == 185 {
			if file.truefilename == file.filename {
			file.truefilename = tcc_strdup(file.filename)
			}
			pstrcpy(file.filename, sizeof(file.filename), &i8(tokc.str.data))
		}
		else if parse_flags & 8 {
		
		}
		else { // 3
		goto _line_err // id: 0x7fffc1b2d3a8
		
}
		n --$
	}
	if file.fd > 0 {
	total_lines += file.line_num - n
	}
	file.line_num = n
	if s1.do_debug {
	put_stabs(file.filename, __stab_debug_code.n_bincl, 0, 0, 0)
	}
	
	}
	 .tok_error, .tok_warning{
	c = tok
	ch = file.buf_ptr [0] 
	skip_spaces()
	q = buf
	for ch != `\n` && ch != (-1) {
		if (q - buf) < sizeof(buf) - 1 {
		*q ++ = ch
		}
		if ch == `\\` {
			if handle_stray_noerror() == 0 {
			q --$
			}
		}
		else { // 3
		inp()
}
	}
	*q = ` `
	if c == Tcc_token.tok_error {
	tcc_error(c'#error %s', buf)
	}
	else { // 3
	tcc_warning(c'#warning %s', buf)
}
	
	}
	 .tok_pragma{ // case comp body kind=CallExpr is_enum=true
	pragma_parse(s1)
	
	}
	 10{ // case comp body kind=GotoStmt is_enum=true
	goto _GOTO_PLACEHOLDER_0x7fffc1b28330 // id: 0x7fffc1b28330
	if tok == `!` && is_bof {
	goto ignore // id: 0x7fffc1b2f110
	}
	tcc_warning(c'Ignoring unknown preprocessing directive #%s', get_tok_str(tok, &tokc))
	// RRRREG ignore id=0x7fffc1b2f110
	ignore: 
	file.buf_ptr = parse_line_comment(file.buf_ptr - 1)
	goto _GOTO_PLACEHOLDER_0x7fffc1b28330 // id: 0x7fffc1b28330
	}
	else {
	if saved_parse_flags & 8 {
	goto ignore // id: 0x7fffc1b2f110
	}
	}
	}
	for tok != 10 {
	next_nomacro()
	}
	// RRRREG the_end id=0x7fffc1b28330
	the_end: 
	parse_flags = saved_parse_flags
}

[export:'ab_month_name']
const (
ab_month_name   = [c'Jan', c'Feb', c'Mar', c'Apr', c'May', c'Jun', c'Jul', c'Aug', c'Sep', c'Oct', c'Nov', c'Dec']!

)

fn next()  {
	if tcc_state.do_debug {
	tcc_debug_line(tcc_state)
	}
	// RRRREG redo id=0x7fffc1b70170
	redo: 
	if parse_flags & 16 {
	next_nomacro_spc()
	}
	else { // 3
	next_nomacro()
}
	if macro_ptr {
		if tok == 204 || tok == 203 {
			goto _GOTO_PLACEHOLDER_0x7fffc1b70170 // id: 0x7fffc1b70170
		}
		else if tok == 0 {
			end_macro()
			goto _GOTO_PLACEHOLDER_0x7fffc1b70170 // id: 0x7fffc1b70170
		}
	}
	else if tok >= 256 && (parse_flags & 1) {
		s := &Sym(0)
		s = define_find(tok)
		if s {
			nested_list := (voidptr(0))
			tokstr_buf.len = 0
			macro_subst_tok(&tokstr_buf, &nested_list, s)
			tok_str_add(&tokstr_buf, 0)
			begin_macro(&tokstr_buf, 0)
			goto _GOTO_PLACEHOLDER_0x7fffc1b70170 // id: 0x7fffc1b70170
		}
	}
	if tok == 190 {
		if parse_flags & 2 {
		parse_number(&i8(tokc.str.data))
		}
	}
	else if tok == 191 {
		if parse_flags & 64 {
		parse_string(&i8(tokc.str.data), tokc.str.size - 1)
		}
	}
}

// skipping global dup "ind"
// skipping global dup "loc"
struct Switch_t { 
	p &&Case_t
	n int
	def_sym int
	bsym &int
	scope &Scope
}
struct Temp_local_variable { 
	location int
	size i16
	align i16
}
struct Scope { 
	prev &Scope
	vla  struct {	loc int
	num int
}

	cl  struct {	s &Sym
	n int
}

	bsym &int
	csym &int
	lstk &Sym
	llstk &Sym
}
fn decl(l int) 

fn gv(rc int) int {
	r := 0
	bit_pos := 0
	bit_size := 0
	size := 0
	align := 0
	rc2 := 0
	
	if vtop.type_.t & 128 {
		type_ := CType{}
		bit_pos = (((vtop.type_.t) >> 20) & 63)
		bit_size = (((vtop.type_.t) >> (20 + 6)) & 63)
		vtop.type_.t &= ~(((1 << (6 + 6)) - 1) << 20 | 128)
		type_.ref = (voidptr(0))
		type_.t = vtop.type_.t & 16
		if (vtop.type_.t & 15) == 11 {
		type_.t |= 16
		}
		r = adjust_bf(vtop, bit_pos, bit_size)
		if (vtop.type_.t & 15) == 4 {
		type_.t |= 4
		}
		else { // 3
		type_.t |= 3
}
		if r == 7 {
			load_packed_bf(&type_, bit_pos, bit_size)
		}
		else {
			bits := if (type_.t & 15) == 4{ 64 } else {32}
			gen_cast(&type_)
			vpushi(bits - (bit_pos + bit_size))
			gen_op(1)
			vpushi(bits - bit_size)
			gen_op(2)
		}
		r = gv(rc)
	}
	else {
		if is_float(vtop.type_.t) && (vtop.r & (63 | 256)) == 48 {
			offset := u32(0)
			size = type_size(&vtop.type_, &align)
			if (nocode_wanted > 0) {
			size = 0 , 1
			align = size = 0
			}
			offset = section_add(data_section, size, align)
			vpush_ref(&vtop.type_, data_section, offset, size)
			vswap()
			init_putv(&vtop.type_, data_section, offset)
			vtop.r |= 256
		}
		if vtop.r & 2048 {
		gbound()
		}
		r = vtop.r & 63
		rc2 = if (rc & 2){ 2 } else {1}
		if rc == 4 {
		rc2 = 16
		}
		else if rc == 4096 {
		rc2 = 8192
		}
		if r >= 48 || (vtop.r & 256) || !(reg_classes [r]  & rc) || ((vtop.type_.t & 15) == 13 && !(reg_classes [vtop.r2]  & rc2)) || ((vtop.type_.t & 15) == 14 && !(reg_classes [vtop.r2]  & rc2)) {
			r = get_reg(rc)
			if ((vtop.type_.t & 15) == 13) || ((vtop.type_.t & 15) == 14) {
				addr_type := 4
load_size := 8
load_type := if ((vtop.type_.t & 15) == 13){ 4 } else {9}

				r2 := 0
				original_type := 0
				
				original_type = vtop.type_.t
				if vtop.r & 256 {
					save_reg_upstack(vtop.r, 1)
					vtop.type_.t = load_type
					load(r, vtop)
					vdup()
					vtop [-1] .r = r
					vtop.type_.t = addr_type
					gaddrof()
					vpushi(load_size)
					gen_op(`+`)
					vtop.r |= 256
					vtop.type_.t = load_type
				}
				else {
					load(r, vtop)
					vdup()
					vtop [-1] .r = r
					vtop.r = vtop [-1] .r2
				}
				r2 = get_reg(rc2)
				load(r2, vtop)
				vpop()
				vtop.r2 = r2
				vtop.type_.t = original_type
			}
			else if (vtop.r & 256) && !is_float(vtop.type_.t) {
				t1 := 0
				t := 0
				
				t = vtop.type_.t
				t1 = t
				if vtop.r & 4096 {
				t = 1
				}
				else if vtop.r & 8192 {
				t = 2
				}
				if vtop.r & 16384 {
				t |= 16
				}
				vtop.type_.t = t
				load(r, vtop)
				vtop.type_.t = t1
			}
			else {
				if vtop.r == 51 {
				vset_vt_jmp()
				}
				load(r, vtop)
			}
		}
		vtop.r = r
	}
	return r
}

fn inc(post int, c int)  {
	test_lvalue()
	vdup()
	if post {
		gv_dup()
		vrotb(3)
		vrotb(3)
	}
	vpushi(c - 163)
	gen_op(`+`)
	vstore()
	if post {
	vpop()
	}
}

fn decl(l int)  {
	decl0(l, 0, (voidptr(0)))
}

struct Dyn_inf { 
	dynamic &Section
	dynstr &Section
	data_offset u32
	rel_addr Elf64_Addr
	rel_size Elf64_Addr
}
fn tcc_output_file(s &TCCState, filename &i8) int {
	ret := 0
	ret = elf_output_file(s, filename)
	return ret
}

struct SectionMergeInfo { 
	s &Section
	offset u32
	new_section u8
	link_once u8
}
struct ArchiveHeader { 
	ar_name [16]i8
	ar_date [12]i8
	ar_uid [6]i8
	ar_gid [6]i8
	ar_mode [8]i8
	ar_size [10]i8
	ar_fmag [2]i8
}
type Sig_t = Sighandler_t
fn tcc_run(s1 &TCCState, argc int, argv &&u8) int {
	prog_main := fn (int, &&i8) int{}
	s1.runtime_main = if s1.nostdlib{ c'_start' } else {c'main'}
	if (s1.dflag & 16) && !find_elf_sym(s1.symtab, s1.runtime_main) {
	return 0
	}
	if tcc_relocate(s1, voidptr(1)) < 0 {
	return -1
	}
	prog_main = tcc_get_symbol_err(s1, s1.runtime_main)
	if s1.do_debug {
		set_exception_handler()
		rt_prog_main = prog_main
	}
	(*__errno_location()) = 0
	if s1.do_bounds_check {
		bound_init := fn (){}
		bound_exit := fn (){}
		bound_new_region := fn (voidptr, Elf64_Addr){}
		bound_delete_region := fn (voidptr) int{}
		i := 0
		ret := 0
		
		rt_bound_error_msg = tcc_get_symbol_err(s1, c'__bound_error_msg')
		bound_init = tcc_get_symbol_err(s1, c'__bound_init')
		bound_exit = tcc_get_symbol_err(s1, c'__bound_exit')
		bound_new_region = tcc_get_symbol_err(s1, c'__bound_new_region')
		bound_delete_region = tcc_get_symbol_err(s1, c'__bound_delete_region')
		bound_init()
		bound_new_region(argv, argc * sizeof(argv [0] ))
		for i = 0 ; i < argc ; i ++ {
		bound_new_region(argv [i] , C.strlen(argv [i] ) + 1)
		}
		ret = (*prog_main)(argc, argv)
		for i = 0 ; i < argc ; i ++ {
		bound_delete_region(argv [i] )
		}
		bound_delete_region(argv)
		bound_exit()
		return ret
	}
	return (*prog_main)(argc, argv)
}

[export:'reg_classes']
const (
reg_classes   = [1 | 4, 1 | 8, 1 | 16, 0, 0, 0, 0, 0, 256, 512, 1024, 2048, 0, 0, 0, 0, 2 | 4096, 2 | 8192, 2 | 16384, 2 | 32768, 2 | 65536, 2 | 131072, 262144, 524288, 128]!

)

fn g(c int)  {
	ind1 := 0
	if nocode_wanted {
	return 
	}
	ind1 = ind + 1
	if ind1 > cur_text_section.data_allocated {
	section_realloc(cur_text_section, ind1)
	}
	cur_text_section.data [ind]  = c
	ind = ind1
}

fn o(c u32)  {
	for c {
		g(c)
		c = c >> 8
	}
}

fn oad(c int, s int) int {
	t := 0
	if nocode_wanted {
	return s
	}
	o(c)
	t = ind
	gen_le32(s)
	return t
}

fn load(r int, sv &SValue)  {
	v := 0
	t := 0
	ft := 0
	fc := 0
	fr := 0
	
	v1 := SValue{}
	fr = sv.r
	ft = sv.type_.t & ~32
	fc = sv..c.i
	if fc != sv..c.i && (fr & 512) {
	tcc_error(c'64 bit addend in load')
	}
	ft &= ~(512 | 256)
	if (fr & 63) == 48 && (fr & 512) && (fr & 256) && !(sv..sym.type_.t & 8192) {
		tr := r | treg_mem
		if is_float(ft) {
			tr = get_reg(1) | treg_mem
		}
		gen_modrm64(139, tr, fr, sv..sym, 0)
		fr = tr | 256
	}
	v = fr & 63
	if fr & 256 {
		b := 0
		ll := 0
		
		if v == 49 {
			v1.type_.t = 5
			v1.r = 50 | 256
			v1..c.i = fc
			fr = r
			if !(reg_classes [fr]  & (1 | 2048)) {
			fr = get_reg(1)
			}
			load(fr, &v1)
		}
		if fc != sv..c.i {
			v1.type_.t = 4
			v1.r = 48
			v1..c.i = sv..c.i
			fr = r
			if !(reg_classes [fr]  & (1 | 2048)) {
			fr = get_reg(1)
			}
			load(fr, &v1)
			fc = 0
		}
		ll = 0
		if (ft & 15) == 7 {
			align := 0
			match type_size(&sv.type_, &align) {
			 1{ // case comp body kind=BinaryOperator is_enum=true
			ft = 1
			
			}
			 2{ // case comp body kind=BinaryOperator is_enum=true
			ft = 2
			
			}
			 4{ // case comp body kind=BinaryOperator is_enum=true
			ft = 3
			
			}
			 8{ // case comp body kind=BinaryOperator is_enum=true
			ft = 4
			
			
			}
			else {
			tcc_error(c'invalid aggregate type for register load')
			}
			}
		}
		if (ft & 15) == 8 {
			b = 7212902
			r = ((r) & 7)
		}
		else if (ft & 15) == 9 {
			b = 8261619
			r = ((r) & 7)
		}
		else if (ft & 15) == 10 {
			b = 219 , 5
			r = b = 219
		}
		else if (ft & (~((4096 | 8192 | 16384 | 32768) | (((1 << (6 + 6)) - 1) << 20 | 128)))) == 1 || (ft & (~((4096 | 8192 | 16384 | 32768) | (((1 << (6 + 6)) - 1) << 20 | 128)))) == 11 {
			b = 48655
		}
		else if (ft & (~((4096 | 8192 | 16384 | 32768) | (((1 << (6 + 6)) - 1) << 20 | 128)))) == (1 | 16) {
			b = 46607
		}
		else if (ft & (~((4096 | 8192 | 16384 | 32768) | (((1 << (6 + 6)) - 1) << 20 | 128)))) == 2 {
			b = 48911
		}
		else if (ft & (~((4096 | 8192 | 16384 | 32768) | (((1 << (6 + 6)) - 1) << 20 | 128)))) == (2 | 16) {
			b = 46863
		}
		else {
			(void(sizeof(if (((ft & 15) == 3) || ((ft & 15) == 4) || ((ft & 15) == 5) || ((ft & 15) == 6)){ 1 } else {0})) , )
			ll = is64_type(ft)
			b = 139
		}
		if ll {
			gen_modrm64(b, r, fr, sv..sym, fc)
		}
		else {
			orex(ll, fr, r, b)
			gen_modrm(r, fr, sv..sym, fc)
		}
	}
	else {
		if v == 48 {
			if fr & 512 {
				if sv..sym.type_.t & 8192 {
					orex(1, 0, r, 141)
					o(5 + ((r) & 7) * 8)
					gen_addrpc32(fr, sv..sym, fc)
				}
				else {
					orex(1, 0, r, 139)
					o(5 + ((r) & 7) * 8)
					gen_gotpcrel(r, sv..sym, fc)
				}
			}
			else if is64_type(ft) {
				orex(1, r, 0, 184 + ((r) & 7))
				gen_le64(sv..c.i)
			}
			else {
				orex(0, r, 0, 184 + ((r) & 7))
				gen_le32(fc)
			}
		}
		else if v == 50 {
			orex(1, 0, r, 141)
			gen_modrm(r, 50, sv..sym, fc)
		}
		else if v == 51 {
			if fc & 256 {
				v = vtop...cmp_r
				fc &= ~256
				orex(0, r, 0, 176 + ((r) & 7))
				g(v ^ fc ^ (v == 149))
				o(890 + ((((r) >> 3) & 1) << 8))
			}
			orex(0, r, 0, 15)
			o(fc)
			o(192 + ((r) & 7))
			orex(0, r, 0, 15)
			o(49334 + ((r) & 7) * 2304)
		}
		else if v == 52 || v == 53 {
			t = v & 1
			orex(0, r, 0, 0)
			oad(184 + ((r) & 7), t)
			o(1515 + ((((r) >> 3) & 1) << 8))
			gsym(fc)
			orex(0, r, 0, 0)
			oad(184 + ((r) & 7), t ^ 1)
		}
		else if v != r {
			if (r >= treg_xmm0) && (r <= treg_xmm7) {
				if v == treg_st0 {
					o(4028914909)
					o(1052658)
					o(68 + ((r) & 7) * 8)
					o(61476)
				}
				else {
					(void(sizeof(if ((v >= treg_xmm0) && (v <= treg_xmm7)){ 1 } else {0})) , )
					if (ft & 15) == 8 {
						o(1052659)
					}
					else {
						(void(sizeof(if ((ft & 15) == 9){ 1 } else {0})) , )
						o(1052658)
					}
					o(192 + ((v) & 7) + ((r) & 7) * 8)
				}
			}
			else if r == treg_st0 {
				(void(sizeof(if ((v >= treg_xmm0) && (v <= treg_xmm7)){ 1 } else {0})) , )
				o(1118194)
				o(68 + ((r) & 7) * 8)
				o(61476)
				o(4028908765)
			}
			else {
				orex(1, r, v, 137)
				o(192 + ((r) & 7) + ((v) & 7) * 8)
			}
		}
	}
}

enum X86_64_Mode {
	x86_64_mode_none
	x86_64_mode_memory
	x86_64_mode_integer
	x86_64_mode_sse
	x86_64_mode_x87
}

[export:'arg_regs']
const (
arg_regs   = [treg_rdi, treg_rsi, treg_rdx, treg_rcx, treg_r8, treg_r9]!

)


const ( // empty enum
	opt_reg8 = 0
	opt_reg16 = 1
	opt_reg32 = 2
	opt_reg64 = 3
	opt_mmx = 4
	opt_sse = 5
	opt_cr = 6
	opt_tr = 7
	opt_db = 8
	opt_seg = 9
	opt_st = 10
	opt_reg8_low = 11
	opt_im8 = 12
	opt_im8s = 13
	opt_im16 = 14
	opt_im32 = 15
	opt_im64 = 16
	opt_eax = 17
	opt_st0 = 18
	opt_cl = 19
	opt_dx = 20
	opt_addr = 21
	opt_indir = 22
	opt_composite_first = 23
	opt_im = 24
	opt_reg = 25
	opt_regw = 26
	opt_imw = 27
	opt_mmxsse = 28
	opt_disp = 29
	opt_disp8 = 30
	opt_ea = 128
)

struct ASMInstr { 
	sym u16
	opcode u16
	instr_type u16
	nb_ops u8
	op_type [3]u8
}
struct Operand { 
	type_ u32
	reg Int8_t
	reg2 Int8_t
	shift u8
	e ExprValue
}
[export:'reg_to_size']
const (
reg_to_size   = [0, 0, 1, 0, 2, 0, 0, 0, 3]!

)

[export:'test_bits']
const (
test_bits   = [0, 1, 2, 2, 2, 3, 3, 3, 4, 4, 5, 5, 6, 6, 7, 7, 8, 9, 10, 10, 11, 11, 12, 12, 13, 13, 14, 14, 15, 15]!

)

[export:'segment_prefixes']
const (
segment_prefixes   = [38, 46, 54, 62, 100, 101]!

)

[export:'asm_instrs']
const (
asm_instrs   = [ASMInstr {
sym: Tcc_token.tok_asm_cmpsb, 
opcode: (u64((if (((166) & 65280) == 3840){ ((((166) >> 8) & ~255) | ((166) & 255)) } else {(166)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((166) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_scmpb, 
opcode: (u64((if (((166) & 65280) == 3840){ ((((166) >> 8) & ~255) | ((166) & 255)) } else {(166)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((166) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_insb, 
opcode: (u64((if (((108) & 65280) == 3840){ ((((108) >> 8) & ~255) | ((108) & 255)) } else {(108)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((108) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_outsb, 
opcode: (u64((if (((110) & 65280) == 3840){ ((((110) >> 8) & ~255) | ((110) & 255)) } else {(110)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((110) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lodsb, 
opcode: (u64((if (((172) & 65280) == 3840){ ((((172) >> 8) & ~255) | ((172) & 255)) } else {(172)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((172) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_slodb, 
opcode: (u64((if (((172) & 65280) == 3840){ ((((172) >> 8) & ~255) | ((172) & 255)) } else {(172)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((172) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movsb, 
opcode: (u64((if (((164) & 65280) == 3840){ ((((164) >> 8) & ~255) | ((164) & 255)) } else {(164)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((164) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_smovb, 
opcode: (u64((if (((164) & 65280) == 3840){ ((((164) >> 8) & ~255) | ((164) & 255)) } else {(164)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((164) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_scasb, 
opcode: (u64((if (((174) & 65280) == 3840){ ((((174) >> 8) & ~255) | ((174) & 255)) } else {(174)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((174) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sscab, 
opcode: (u64((if (((174) & 65280) == 3840){ ((((174) >> 8) & ~255) | ((174) & 255)) } else {(174)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((174) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_stosb, 
opcode: (u64((if (((170) & 65280) == 3840){ ((((170) >> 8) & ~255) | ((170) & 255)) } else {(170)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((170) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sstob, 
opcode: (u64((if (((170) & 65280) == 3840){ ((((170) >> 8) & ~255) | ((170) & 255)) } else {(170)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((170) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_bsfw, 
opcode: (u64((if (((4028) & 65280) == 3840){ ((((4028) >> 8) & ~255) | ((4028) & 255)) } else {(4028)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4028) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_bsrw, 
opcode: (u64((if (((4029) & 65280) == 3840){ ((((4029) >> 8) & ~255) | ((4029) & 255)) } else {(4029)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4029) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btw, 
opcode: (u64((if (((4003) & 65280) == 3840){ ((((4003) >> 8) & ~255) | ((4003) & 255)) } else {(4003)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4003) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btw, 
opcode: (u64((if (((4026) & 65280) == 3840){ ((((4026) >> 8) & ~255) | ((4026) & 255)) } else {(4026)}))), 
instr_type: ((8 | 4096) | ((4) << 13) | (if (((4026) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btsw, 
opcode: (u64((if (((4011) & 65280) == 3840){ ((((4011) >> 8) & ~255) | ((4011) & 255)) } else {(4011)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4011) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btsw, 
opcode: (u64((if (((4026) & 65280) == 3840){ ((((4026) >> 8) & ~255) | ((4026) & 255)) } else {(4026)}))), 
instr_type: ((8 | 4096) | ((5) << 13) | (if (((4026) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btrw, 
opcode: (u64((if (((4019) & 65280) == 3840){ ((((4019) >> 8) & ~255) | ((4019) & 255)) } else {(4019)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4019) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btrw, 
opcode: (u64((if (((4026) & 65280) == 3840){ ((((4026) >> 8) & ~255) | ((4026) & 255)) } else {(4026)}))), 
instr_type: ((8 | 4096) | ((6) << 13) | (if (((4026) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btcw, 
opcode: (u64((if (((4027) & 65280) == 3840){ ((((4027) >> 8) & ~255) | ((4027) & 255)) } else {(4027)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4027) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_btcw, 
opcode: (u64((if (((4026) & 65280) == 3840){ ((((4026) >> 8) & ~255) | ((4026) & 255)) } else {(4026)}))), 
instr_type: ((8 | 4096) | ((7) << 13) | (if (((4026) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sysretq, 
opcode: (u64((if (((4722439) & 65280) == 3840){ ((((4722439) >> 8) & ~255) | ((4722439) & 255)) } else {(4722439)}))), 
instr_type: ((0) | ((0) << 13) | (if (((4722439) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movb, 
opcode: (u64((if (((136) & 65280) == 3840){ ((((136) >> 8) & ~255) | ((136) & 255)) } else {(136)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((136) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movb, 
opcode: (u64((if (((138) & 65280) == 3840){ ((((138) >> 8) & ~255) | ((138) & 255)) } else {(138)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((138) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movb, 
opcode: (u64((if (((176) & 65280) == 3840){ ((((176) >> 8) & ~255) | ((176) & 255)) } else {(176)}))), 
instr_type: ((4 | (1 | 4096)) | ((0) << 13) | (if (((176) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_mov, 
opcode: (u64((if (((184) & 65280) == 3840){ ((((184) >> 8) & ~255) | ((184) & 255)) } else {(184)}))), 
instr_type: ((4) | ((0) << 13) | (if (((184) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im64, opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((184) & 65280) == 3840){ ((((184) >> 8) & ~255) | ((184) & 255)) } else {(184)}))), 
instr_type: ((4) | ((0) << 13) | (if (((184) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im64, opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movb, 
opcode: (u64((if (((198) & 65280) == 3840){ ((((198) >> 8) & ~255) | ((198) & 255)) } else {(198)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((198) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((140) & 65280) == 3840){ ((((140) >> 8) & ~255) | ((140) & 255)) } else {(140)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((140) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_seg, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((142) & 65280) == 3840){ ((((142) >> 8) & ~255) | ((142) & 255)) } else {(142)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((142) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_seg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((3872) & 65280) == 3840){ ((((3872) >> 8) & ~255) | ((3872) & 255)) } else {(3872)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3872) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_cr, opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((3873) & 65280) == 3840){ ((((3873) >> 8) & ~255) | ((3873) & 255)) } else {(3873)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3873) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_db, opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((3874) & 65280) == 3840){ ((((3874) >> 8) & ~255) | ((3874) & 255)) } else {(3874)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3874) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg64, opt_cr]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movw, 
opcode: (u64((if (((3875) & 65280) == 3840){ ((((3875) >> 8) & ~255) | ((3875) & 255)) } else {(3875)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3875) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg64, opt_db]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movsbw, 
opcode: (u64((if (((6688702) & 65280) == 3840){ ((((6688702) >> 8) & ~255) | ((6688702) & 255)) } else {(6688702)}))), 
instr_type: ((8) | ((0) << 13) | (if (((6688702) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg8 | opt_ea, opt_reg16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movsbl, 
opcode: (u64((if (((4030) & 65280) == 3840){ ((((4030) >> 8) & ~255) | ((4030) & 255)) } else {(4030)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4030) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg8 | opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movsbq, 
opcode: (u64((if (((4030) & 65280) == 3840){ ((((4030) >> 8) & ~255) | ((4030) & 255)) } else {(4030)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4030) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg8 | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movswl, 
opcode: (u64((if (((4031) & 65280) == 3840){ ((((4031) >> 8) & ~255) | ((4031) & 255)) } else {(4031)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4031) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg16 | opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movswq, 
opcode: (u64((if (((4031) & 65280) == 3840){ ((((4031) >> 8) & ~255) | ((4031) & 255)) } else {(4031)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4031) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg16 | opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movslq, 
opcode: (u64((if (((99) & 65280) == 3840){ ((((99) >> 8) & ~255) | ((99) & 255)) } else {(99)}))), 
instr_type: ((8) | ((0) << 13) | (if (((99) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg32 | opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movzbw, 
opcode: (u64((if (((4022) & 65280) == 3840){ ((((4022) >> 8) & ~255) | ((4022) & 255)) } else {(4022)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4022) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg8 | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movzwl, 
opcode: (u64((if (((4023) & 65280) == 3840){ ((((4023) >> 8) & ~255) | ((4023) & 255)) } else {(4023)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4023) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg16 | opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movzwq, 
opcode: (u64((if (((4023) & 65280) == 3840){ ((((4023) >> 8) & ~255) | ((4023) & 255)) } else {(4023)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4023) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg16 | opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushq, 
opcode: (u64((if (((106) & 65280) == 3840){ ((((106) >> 8) & ~255) | ((106) & 255)) } else {(106)}))), 
instr_type: ((0) | ((0) << 13) | (if (((106) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8s]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_push, 
opcode: (u64((if (((106) & 65280) == 3840){ ((((106) >> 8) & ~255) | ((106) & 255)) } else {(106)}))), 
instr_type: ((0) | ((0) << 13) | (if (((106) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8s]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((26218) & 65280) == 3840){ ((((26218) >> 8) & ~255) | ((26218) & 255)) } else {(26218)}))), 
instr_type: ((0) | ((0) << 13) | (if (((26218) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8s]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((80) & 65280) == 3840){ ((((80) >> 8) & ~255) | ((80) & 255)) } else {(80)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((80) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((80) & 65280) == 3840){ ((((80) >> 8) & ~255) | ((80) & 255)) } else {(80)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((80) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8 | 4096) | ((6) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg64 | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((26216) & 65280) == 3840){ ((((26216) >> 8) & ~255) | ((26216) & 255)) } else {(26216)}))), 
instr_type: ((0) | ((0) << 13) | (if (((26216) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((104) & 65280) == 3840){ ((((104) >> 8) & ~255) | ((104) & 255)) } else {(104)}))), 
instr_type: ((4096) | ((0) << 13) | (if (((104) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pushw, 
opcode: (u64((if (((6) & 65280) == 3840){ ((((6) >> 8) & ~255) | ((6) & 255)) } else {(6)}))), 
instr_type: ((4096) | ((0) << 13) | (if (((6) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_seg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_popw, 
opcode: (u64((if (((88) & 65280) == 3840){ ((((88) >> 8) & ~255) | ((88) & 255)) } else {(88)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((88) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_popw, 
opcode: (u64((if (((88) & 65280) == 3840){ ((((88) >> 8) & ~255) | ((88) & 255)) } else {(88)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((88) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_popw, 
opcode: (u64((if (((143) & 65280) == 3840){ ((((143) >> 8) & ~255) | ((143) & 255)) } else {(143)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((143) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_regw | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_popw, 
opcode: (u64((if (((7) & 65280) == 3840){ ((((7) >> 8) & ~255) | ((7) & 255)) } else {(7)}))), 
instr_type: ((4096) | ((0) << 13) | (if (((7) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_seg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_xchgw, 
opcode: (u64((if (((144) & 65280) == 3840){ ((((144) >> 8) & ~255) | ((144) & 255)) } else {(144)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((144) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_xchgw, 
opcode: (u64((if (((144) & 65280) == 3840){ ((((144) >> 8) & ~255) | ((144) & 255)) } else {(144)}))), 
instr_type: ((4 | 4096) | ((0) << 13) | (if (((144) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_eax, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_xchgb, 
opcode: (u64((if (((134) & 65280) == 3840){ ((((134) >> 8) & ~255) | ((134) & 255)) } else {(134)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((134) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_xchgb, 
opcode: (u64((if (((134) & 65280) == 3840){ ((((134) >> 8) & ~255) | ((134) & 255)) } else {(134)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((134) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_inb, 
opcode: (u64((if (((228) & 65280) == 3840){ ((((228) >> 8) & ~255) | ((228) & 255)) } else {(228)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((228) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_inb, 
opcode: (u64((if (((228) & 65280) == 3840){ ((((228) >> 8) & ~255) | ((228) & 255)) } else {(228)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((228) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_inb, 
opcode: (u64((if (((236) & 65280) == 3840){ ((((236) >> 8) & ~255) | ((236) & 255)) } else {(236)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((236) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_dx, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_inb, 
opcode: (u64((if (((236) & 65280) == 3840){ ((((236) >> 8) & ~255) | ((236) & 255)) } else {(236)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((236) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_dx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_outb, 
opcode: (u64((if (((230) & 65280) == 3840){ ((((230) >> 8) & ~255) | ((230) & 255)) } else {(230)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((230) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_eax, opt_im8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_outb, 
opcode: (u64((if (((230) & 65280) == 3840){ ((((230) >> 8) & ~255) | ((230) & 255)) } else {(230)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((230) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_outb, 
opcode: (u64((if (((238) & 65280) == 3840){ ((((238) >> 8) & ~255) | ((238) & 255)) } else {(238)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((238) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_eax, opt_dx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_outb, 
opcode: (u64((if (((238) & 65280) == 3840){ ((((238) >> 8) & ~255) | ((238) & 255)) } else {(238)}))), 
instr_type: (((1 | 2)) | ((0) << 13) | (if (((238) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_dx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_leaw, 
opcode: (u64((if (((141) & 65280) == 3840){ ((((141) >> 8) & ~255) | ((141) & 255)) } else {(141)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((141) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_les, 
opcode: (u64((if (((196) & 65280) == 3840){ ((((196) >> 8) & ~255) | ((196) & 255)) } else {(196)}))), 
instr_type: ((8) | ((0) << 13) | (if (((196) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lds, 
opcode: (u64((if (((197) & 65280) == 3840){ ((((197) >> 8) & ~255) | ((197) & 255)) } else {(197)}))), 
instr_type: ((8) | ((0) << 13) | (if (((197) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lss, 
opcode: (u64((if (((4018) & 65280) == 3840){ ((((4018) >> 8) & ~255) | ((4018) & 255)) } else {(4018)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4018) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lfs, 
opcode: (u64((if (((4020) & 65280) == 3840){ ((((4020) >> 8) & ~255) | ((4020) & 255)) } else {(4020)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4020) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lgs, 
opcode: (u64((if (((4021) & 65280) == 3840){ ((((4021) >> 8) & ~255) | ((4021) & 255)) } else {(4021)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4021) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea, opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addb, 
opcode: (u64((if (((0) & 65280) == 3840){ ((((0) >> 8) & ~255) | ((0) & 255)) } else {(0)}))), 
instr_type: ((48 | 8 | (1 | 4096)) | ((0) << 13) | (if (((0) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addb, 
opcode: (u64((if (((2) & 65280) == 3840){ ((((2) >> 8) & ~255) | ((2) & 255)) } else {(2)}))), 
instr_type: ((48 | 8 | (1 | 4096)) | ((0) << 13) | (if (((2) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addb, 
opcode: (u64((if (((4) & 65280) == 3840){ ((((4) >> 8) & ~255) | ((4) & 255)) } else {(4)}))), 
instr_type: ((48 | (1 | 4096)) | ((0) << 13) | (if (((4) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addw, 
opcode: (u64((if (((131) & 65280) == 3840){ ((((131) >> 8) & ~255) | ((131) & 255)) } else {(131)}))), 
instr_type: ((48 | 8 | 4096) | ((0) << 13) | (if (((131) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8s, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addb, 
opcode: (u64((if (((128) & 65280) == 3840){ ((((128) >> 8) & ~255) | ((128) & 255)) } else {(128)}))), 
instr_type: ((48 | 8 | (1 | 4096)) | ((0) << 13) | (if (((128) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_testb, 
opcode: (u64((if (((132) & 65280) == 3840){ ((((132) >> 8) & ~255) | ((132) & 255)) } else {(132)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((132) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_testb, 
opcode: (u64((if (((132) & 65280) == 3840){ ((((132) >> 8) & ~255) | ((132) & 255)) } else {(132)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((132) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_testb, 
opcode: (u64((if (((168) & 65280) == 3840){ ((((168) >> 8) & ~255) | ((168) & 255)) } else {(168)}))), 
instr_type: (((1 | 4096)) | ((0) << 13) | (if (((168) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_testb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_incb, 
opcode: (u64((if (((254) & 65280) == 3840){ ((((254) >> 8) & ~255) | ((254) & 255)) } else {(254)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((254) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_decb, 
opcode: (u64((if (((254) & 65280) == 3840){ ((((254) >> 8) & ~255) | ((254) & 255)) } else {(254)}))), 
instr_type: ((8 | (1 | 4096)) | ((1) << 13) | (if (((254) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_notb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((2) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_negb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((3) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_mulb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((4) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((5) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulw, 
opcode: (u64((if (((4015) & 65280) == 3840){ ((((4015) >> 8) & ~255) | ((4015) & 255)) } else {(4015)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4015) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg | opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulw, 
opcode: (u64((if (((107) & 65280) == 3840){ ((((107) >> 8) & ~255) | ((107) & 255)) } else {(107)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((107) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_im8s, opt_regw | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulw, 
opcode: (u64((if (((107) & 65280) == 3840){ ((((107) >> 8) & ~255) | ((107) & 255)) } else {(107)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((107) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8s, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulw, 
opcode: (u64((if (((105) & 65280) == 3840){ ((((105) >> 8) & ~255) | ((105) & 255)) } else {(105)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((105) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_imw, opt_regw | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_imulw, 
opcode: (u64((if (((105) & 65280) == 3840){ ((((105) >> 8) & ~255) | ((105) & 255)) } else {(105)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((105) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_imw, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_divb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((6) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_divb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((6) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg | opt_ea, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_idivb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((7) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_idivb, 
opcode: (u64((if (((246) & 65280) == 3840){ ((((246) >> 8) & ~255) | ((246) & 255)) } else {(246)}))), 
instr_type: ((8 | (1 | 4096)) | ((7) << 13) | (if (((246) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg | opt_ea, opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_rolb, 
opcode: (u64((if (((192) & 65280) == 3840){ ((((192) >> 8) & ~255) | ((192) & 255)) } else {(192)}))), 
instr_type: ((8 | (1 | 4096) | 32) | ((0) << 13) | (if (((192) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_rolb, 
opcode: (u64((if (((210) & 65280) == 3840){ ((((210) >> 8) & ~255) | ((210) & 255)) } else {(210)}))), 
instr_type: ((8 | (1 | 4096) | 32) | ((0) << 13) | (if (((210) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_cl, opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_rolb, 
opcode: (u64((if (((208) & 65280) == 3840){ ((((208) >> 8) & ~255) | ((208) & 255)) } else {(208)}))), 
instr_type: ((8 | (1 | 4096) | 32) | ((0) << 13) | (if (((208) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shldw, 
opcode: (u64((if (((4004) & 65280) == 3840){ ((((4004) >> 8) & ~255) | ((4004) & 255)) } else {(4004)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4004) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_im8, opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shldw, 
opcode: (u64((if (((4005) & 65280) == 3840){ ((((4005) >> 8) & ~255) | ((4005) & 255)) } else {(4005)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4005) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_cl, opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shldw, 
opcode: (u64((if (((4005) & 65280) == 3840){ ((((4005) >> 8) & ~255) | ((4005) & 255)) } else {(4005)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4005) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shrdw, 
opcode: (u64((if (((4012) & 65280) == 3840){ ((((4012) >> 8) & ~255) | ((4012) & 255)) } else {(4012)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4012) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_im8, opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shrdw, 
opcode: (u64((if (((4013) & 65280) == 3840){ ((((4013) >> 8) & ~255) | ((4013) & 255)) } else {(4013)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4013) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 3, 
op_type: [opt_cl, opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_shrdw, 
opcode: (u64((if (((4013) & 65280) == 3840){ ((((4013) >> 8) & ~255) | ((4013) & 255)) } else {(4013)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((4013) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw, opt_ea | opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_call, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8) | ((2) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_indir]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_call, 
opcode: (u64((if (((232) & 65280) == 3840){ ((((232) >> 8) & ~255) | ((232) & 255)) } else {(232)}))), 
instr_type: ((0) | ((0) << 13) | (if (((232) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_jmp, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8) | ((4) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_indir]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_jmp, 
opcode: (u64((if (((235) & 65280) == 3840){ ((((235) >> 8) & ~255) | ((235) & 255)) } else {(235)}))), 
instr_type: ((0) | ((0) << 13) | (if (((235) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lcall, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8) | ((3) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ljmp, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8) | ((5) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ljmpw, 
opcode: (u64((if (((26367) & 65280) == 3840){ ((((26367) >> 8) & ~255) | ((26367) & 255)) } else {(26367)}))), 
instr_type: ((8) | ((5) << 13) | (if (((26367) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ljmpl, 
opcode: (u64((if (((255) & 65280) == 3840){ ((((255) >> 8) & ~255) | ((255) & 255)) } else {(255)}))), 
instr_type: ((8) | ((5) << 13) | (if (((255) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_int, 
opcode: (u64((if (((205) & 65280) == 3840){ ((((205) >> 8) & ~255) | ((205) & 255)) } else {(205)}))), 
instr_type: ((0) | ((0) << 13) | (if (((205) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_seto, 
opcode: (u64((if (((3984) & 65280) == 3840){ ((((3984) >> 8) & ~255) | ((3984) & 255)) } else {(3984)}))), 
instr_type: ((8 | 80) | ((0) << 13) | (if (((3984) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg8 | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_setob, 
opcode: (u64((if (((3984) & 65280) == 3840){ ((((3984) >> 8) & ~255) | ((3984) & 255)) } else {(3984)}))), 
instr_type: ((8 | 80) | ((0) << 13) | (if (((3984) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg8 | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_enter, 
opcode: (u64((if (((200) & 65280) == 3840){ ((((200) >> 8) & ~255) | ((200) & 255)) } else {(200)}))), 
instr_type: ((0) | ((0) << 13) | (if (((200) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im16, opt_im8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_retq, 
opcode: (u64((if (((194) & 65280) == 3840){ ((((194) >> 8) & ~255) | ((194) & 255)) } else {(194)}))), 
instr_type: ((0) | ((0) << 13) | (if (((194) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ret, 
opcode: (u64((if (((194) & 65280) == 3840){ ((((194) >> 8) & ~255) | ((194) & 255)) } else {(194)}))), 
instr_type: ((0) | ((0) << 13) | (if (((194) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lret, 
opcode: (u64((if (((202) & 65280) == 3840){ ((((202) >> 8) & ~255) | ((202) & 255)) } else {(202)}))), 
instr_type: ((0) | ((0) << 13) | (if (((202) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_im16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_jo, 
opcode: (u64((if (((112) & 65280) == 3840){ ((((112) >> 8) & ~255) | ((112) & 255)) } else {(112)}))), 
instr_type: ((80) | ((0) << 13) | (if (((112) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_loopne, 
opcode: (u64((if (((224) & 65280) == 3840){ ((((224) >> 8) & ~255) | ((224) & 255)) } else {(224)}))), 
instr_type: ((0) | ((0) << 13) | (if (((224) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_loopnz, 
opcode: (u64((if (((224) & 65280) == 3840){ ((((224) >> 8) & ~255) | ((224) & 255)) } else {(224)}))), 
instr_type: ((0) | ((0) << 13) | (if (((224) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_loope, 
opcode: (u64((if (((225) & 65280) == 3840){ ((((225) >> 8) & ~255) | ((225) & 255)) } else {(225)}))), 
instr_type: ((0) | ((0) << 13) | (if (((225) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_loopz, 
opcode: (u64((if (((225) & 65280) == 3840){ ((((225) >> 8) & ~255) | ((225) & 255)) } else {(225)}))), 
instr_type: ((0) | ((0) << 13) | (if (((225) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_loop, 
opcode: (u64((if (((226) & 65280) == 3840){ ((((226) >> 8) & ~255) | ((226) & 255)) } else {(226)}))), 
instr_type: ((0) | ((0) << 13) | (if (((226) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_jecxz, 
opcode: (u64((if (((26595) & 65280) == 3840){ ((((26595) >> 8) & ~255) | ((26595) & 255)) } else {(26595)}))), 
instr_type: ((0) | ((0) << 13) | (if (((26595) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_disp8]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcomp, 
opcode: (u64((if (((55513) & 65280) == 3840){ ((((55513) >> 8) & ~255) | ((55513) & 255)) } else {(55513)}))), 
instr_type: ((0) | ((0) << 13) | (if (((55513) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fadd, 
opcode: (u64((if (((55488) & 65280) == 3840){ ((((55488) >> 8) & ~255) | ((55488) & 255)) } else {(55488)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((55488) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fadd, 
opcode: (u64((if (((55488) & 65280) == 3840){ ((((55488) >> 8) & ~255) | ((55488) & 255)) } else {(55488)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((55488) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fadd, 
opcode: (u64((if (((56512) & 65280) == 3840){ ((((56512) >> 8) & ~255) | ((56512) & 255)) } else {(56512)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((56512) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st0, opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fmul, 
opcode: (u64((if (((56520) & 65280) == 3840){ ((((56520) >> 8) & ~255) | ((56520) & 255)) } else {(56520)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((56520) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st0, opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fadd, 
opcode: (u64((if (((57025) & 65280) == 3840){ ((((57025) >> 8) & ~255) | ((57025) & 255)) } else {(57025)}))), 
instr_type: ((64) | ((0) << 13) | (if (((57025) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_faddp, 
opcode: (u64((if (((57024) & 65280) == 3840){ ((((57024) >> 8) & ~255) | ((57024) & 255)) } else {(57024)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((57024) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_faddp, 
opcode: (u64((if (((57024) & 65280) == 3840){ ((((57024) >> 8) & ~255) | ((57024) & 255)) } else {(57024)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((57024) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_faddp, 
opcode: (u64((if (((57024) & 65280) == 3840){ ((((57024) >> 8) & ~255) | ((57024) & 255)) } else {(57024)}))), 
instr_type: ((64 | 4) | ((0) << 13) | (if (((57024) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st0, opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_faddp, 
opcode: (u64((if (((57025) & 65280) == 3840){ ((((57025) >> 8) & ~255) | ((57025) & 255)) } else {(57025)}))), 
instr_type: ((64) | ((0) << 13) | (if (((57025) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fadds, 
opcode: (u64((if (((216) & 65280) == 3840){ ((((216) >> 8) & ~255) | ((216) & 255)) } else {(216)}))), 
instr_type: ((64 | 8) | ((0) << 13) | (if (((216) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fiaddl, 
opcode: (u64((if (((218) & 65280) == 3840){ ((((218) >> 8) & ~255) | ((218) & 255)) } else {(218)}))), 
instr_type: ((64 | 8) | ((0) << 13) | (if (((218) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_faddl, 
opcode: (u64((if (((220) & 65280) == 3840){ ((((220) >> 8) & ~255) | ((220) & 255)) } else {(220)}))), 
instr_type: ((64 | 8) | ((0) << 13) | (if (((220) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fiadds, 
opcode: (u64((if (((222) & 65280) == 3840){ ((((222) >> 8) & ~255) | ((222) & 255)) } else {(222)}))), 
instr_type: ((64 | 8) | ((0) << 13) | (if (((222) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fld, 
opcode: (u64((if (((55744) & 65280) == 3840){ ((((55744) >> 8) & ~255) | ((55744) & 255)) } else {(55744)}))), 
instr_type: ((4) | ((0) << 13) | (if (((55744) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fldl, 
opcode: (u64((if (((55744) & 65280) == 3840){ ((((55744) >> 8) & ~255) | ((55744) & 255)) } else {(55744)}))), 
instr_type: ((4) | ((0) << 13) | (if (((55744) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_flds, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((0) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fldl, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((0) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fildl, 
opcode: (u64((if (((219) & 65280) == 3840){ ((((219) >> 8) & ~255) | ((219) & 255)) } else {(219)}))), 
instr_type: ((8) | ((0) << 13) | (if (((219) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fildq, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((5) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fildll, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((5) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fldt, 
opcode: (u64((if (((219) & 65280) == 3840){ ((((219) >> 8) & ~255) | ((219) & 255)) } else {(219)}))), 
instr_type: ((8) | ((5) << 13) | (if (((219) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fbld, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((4) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fst, 
opcode: (u64((if (((56784) & 65280) == 3840){ ((((56784) >> 8) & ~255) | ((56784) & 255)) } else {(56784)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56784) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstl, 
opcode: (u64((if (((56784) & 65280) == 3840){ ((((56784) >> 8) & ~255) | ((56784) & 255)) } else {(56784)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56784) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fsts, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((2) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstps, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((3) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstl, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((2) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstpl, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((3) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fist, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((2) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fistp, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((3) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fistl, 
opcode: (u64((if (((219) & 65280) == 3840){ ((((219) >> 8) & ~255) | ((219) & 255)) } else {(219)}))), 
instr_type: ((8) | ((2) << 13) | (if (((219) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fistpl, 
opcode: (u64((if (((219) & 65280) == 3840){ ((((219) >> 8) & ~255) | ((219) & 255)) } else {(219)}))), 
instr_type: ((8) | ((3) << 13) | (if (((219) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstp, 
opcode: (u64((if (((56792) & 65280) == 3840){ ((((56792) >> 8) & ~255) | ((56792) & 255)) } else {(56792)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56792) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fistpq, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((7) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fistpll, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((7) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstpt, 
opcode: (u64((if (((219) & 65280) == 3840){ ((((219) >> 8) & ~255) | ((219) & 255)) } else {(219)}))), 
instr_type: ((8) | ((7) << 13) | (if (((219) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fbstp, 
opcode: (u64((if (((223) & 65280) == 3840){ ((((223) >> 8) & ~255) | ((223) & 255)) } else {(223)}))), 
instr_type: ((8) | ((6) << 13) | (if (((223) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fxch, 
opcode: (u64((if (((55752) & 65280) == 3840){ ((((55752) >> 8) & ~255) | ((55752) & 255)) } else {(55752)}))), 
instr_type: ((4) | ((0) << 13) | (if (((55752) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fucom, 
opcode: (u64((if (((56800) & 65280) == 3840){ ((((56800) >> 8) & ~255) | ((56800) & 255)) } else {(56800)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56800) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fucomp, 
opcode: (u64((if (((56808) & 65280) == 3840){ ((((56808) >> 8) & ~255) | ((56808) & 255)) } else {(56808)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56808) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_finit, 
opcode: (u64((if (((56291) & 65280) == 3840){ ((((56291) >> 8) & ~255) | ((56291) & 255)) } else {(56291)}))), 
instr_type: ((16) | ((0) << 13) | (if (((56291) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fldcw, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((5) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fnstcw, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((7) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstcw, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8 | 16) | ((7) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fnstsw, 
opcode: (u64((if (((57312) & 65280) == 3840){ ((((57312) >> 8) & ~255) | ((57312) & 255)) } else {(57312)}))), 
instr_type: ((0) | ((0) << 13) | (if (((57312) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fnstsw, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((7) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstsw, 
opcode: (u64((if (((57312) & 65280) == 3840){ ((((57312) >> 8) & ~255) | ((57312) & 255)) } else {(57312)}))), 
instr_type: ((16) | ((0) << 13) | (if (((57312) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_eax]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstsw, 
opcode: (u64((if (((57312) & 65280) == 3840){ ((((57312) >> 8) & ~255) | ((57312) & 255)) } else {(57312)}))), 
instr_type: ((16) | ((0) << 13) | (if (((57312) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstsw, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8 | 16) | ((7) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fclex, 
opcode: (u64((if (((56290) & 65280) == 3840){ ((((56290) >> 8) & ~255) | ((56290) & 255)) } else {(56290)}))), 
instr_type: ((16) | ((0) << 13) | (if (((56290) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fnstenv, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((6) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fstenv, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8 | 16) | ((6) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fldenv, 
opcode: (u64((if (((217) & 65280) == 3840){ ((((217) >> 8) & ~255) | ((217) & 255)) } else {(217)}))), 
instr_type: ((8) | ((4) << 13) | (if (((217) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fnsave, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((6) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fsave, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8 | 16) | ((6) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_frstor, 
opcode: (u64((if (((221) & 65280) == 3840){ ((((221) >> 8) & ~255) | ((221) & 255)) } else {(221)}))), 
instr_type: ((8) | ((4) << 13) | (if (((221) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ffree, 
opcode: (u64((if (((56768) & 65280) == 3840){ ((((56768) >> 8) & ~255) | ((56768) & 255)) } else {(56768)}))), 
instr_type: ((4) | ((4) << 13) | (if (((56768) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ffreep, 
opcode: (u64((if (((57280) & 65280) == 3840){ ((((57280) >> 8) & ~255) | ((57280) & 255)) } else {(57280)}))), 
instr_type: ((4) | ((4) << 13) | (if (((57280) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_st]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fxsave, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fxrstor, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((1) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fxsaveq, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8 | 512) | ((0) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fxrstorq, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8 | 512) | ((1) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_arpl, 
opcode: (u64((if (((99) & 65280) == 3840){ ((((99) >> 8) & ~255) | ((99) & 255)) } else {(99)}))), 
instr_type: ((8) | ((0) << 13) | (if (((99) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg16, opt_reg16 | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_larw, 
opcode: (u64((if (((3842) & 65280) == 3840){ ((((3842) >> 8) & ~255) | ((3842) & 255)) } else {(3842)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3842) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg | opt_ea, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lgdt, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lgdtq, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lidt, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((3) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lidtq, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((3) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lldt, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lmsw, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((6) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea | opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lslw, 
opcode: (u64((if (((3843) & 65280) == 3840){ ((((3843) >> 8) & ~255) | ((3843) & 255)) } else {(3843)}))), 
instr_type: ((8 | 4096) | ((0) << 13) | (if (((3843) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg, opt_reg]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_ltr, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((3) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea | opt_reg16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sgdt, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sgdtq, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sidt, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((1) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sidtq, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((1) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sldt, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_smsw, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((4) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_str, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((1) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg32 | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_str, 
opcode: (u64((if (((6688512) & 65280) == 3840){ ((((6688512) >> 8) & ~255) | ((6688512) & 255)) } else {(6688512)}))), 
instr_type: ((8) | ((1) << 13) | (if (((6688512) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg16]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_str, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8 | 512) | ((1) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_verr, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((4) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_verw, 
opcode: (u64((if (((3840) & 65280) == 3840){ ((((3840) >> 8) & ~255) | ((3840) & 255)) } else {(3840)}))), 
instr_type: ((8) | ((5) << 13) | (if (((3840) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_swapgs, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((7) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_bswap, 
opcode: (u64((if (((4040) & 65280) == 3840){ ((((4040) >> 8) & ~255) | ((4040) & 255)) } else {(4040)}))), 
instr_type: ((4) | ((0) << 13) | (if (((4040) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_bswapl, 
opcode: (u64((if (((4040) & 65280) == 3840){ ((((4040) >> 8) & ~255) | ((4040) & 255)) } else {(4040)}))), 
instr_type: ((4) | ((0) << 13) | (if (((4040) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_bswapq, 
opcode: (u64((if (((4040) & 65280) == 3840){ ((((4040) >> 8) & ~255) | ((4040) & 255)) } else {(4040)}))), 
instr_type: ((4 | 512) | ((0) << 13) | (if (((4040) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_xaddb, 
opcode: (u64((if (((4032) & 65280) == 3840){ ((((4032) >> 8) & ~255) | ((4032) & 255)) } else {(4032)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((4032) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cmpxchgb, 
opcode: (u64((if (((4016) & 65280) == 3840){ ((((4016) >> 8) & ~255) | ((4016) & 255)) } else {(4016)}))), 
instr_type: ((8 | (1 | 4096)) | ((0) << 13) | (if (((4016) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg, opt_reg | opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_invlpg, 
opcode: (u64((if (((3841) & 65280) == 3840){ ((((3841) >> 8) & ~255) | ((3841) & 255)) } else {(3841)}))), 
instr_type: ((8) | ((7) << 13) | (if (((3841) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cmpxchg8b, 
opcode: (u64((if (((4039) & 65280) == 3840){ ((((4039) >> 8) & ~255) | ((4039) & 255)) } else {(4039)}))), 
instr_type: ((8) | ((1) << 13) | (if (((4039) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cmpxchg16b, 
opcode: (u64((if (((4039) & 65280) == 3840){ ((((4039) >> 8) & ~255) | ((4039) & 255)) } else {(4039)}))), 
instr_type: ((8 | 512) | ((1) << 13) | (if (((4039) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cmovo, 
opcode: (u64((if (((3904) & 65280) == 3840){ ((((3904) >> 8) & ~255) | ((3904) & 255)) } else {(3904)}))), 
instr_type: ((8 | 80 | 4096) | ((0) << 13) | (if (((3904) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_regw | opt_ea, opt_regw]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovb, 
opcode: (u64((if (((56000) & 65280) == 3840){ ((((56000) >> 8) & ~255) | ((56000) & 255)) } else {(56000)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56000) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmove, 
opcode: (u64((if (((56008) & 65280) == 3840){ ((((56008) >> 8) & ~255) | ((56008) & 255)) } else {(56008)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56008) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovbe, 
opcode: (u64((if (((56016) & 65280) == 3840){ ((((56016) >> 8) & ~255) | ((56016) & 255)) } else {(56016)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56016) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovu, 
opcode: (u64((if (((56024) & 65280) == 3840){ ((((56024) >> 8) & ~255) | ((56024) & 255)) } else {(56024)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56024) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovnb, 
opcode: (u64((if (((56256) & 65280) == 3840){ ((((56256) >> 8) & ~255) | ((56256) & 255)) } else {(56256)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56256) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovne, 
opcode: (u64((if (((56264) & 65280) == 3840){ ((((56264) >> 8) & ~255) | ((56264) & 255)) } else {(56264)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56264) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovnbe, 
opcode: (u64((if (((56272) & 65280) == 3840){ ((((56272) >> 8) & ~255) | ((56272) & 255)) } else {(56272)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56272) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcmovnu, 
opcode: (u64((if (((56280) & 65280) == 3840){ ((((56280) >> 8) & ~255) | ((56280) & 255)) } else {(56280)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56280) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fucomi, 
opcode: (u64((if (((56296) & 65280) == 3840){ ((((56296) >> 8) & ~255) | ((56296) & 255)) } else {(56296)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56296) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcomi, 
opcode: (u64((if (((56304) & 65280) == 3840){ ((((56304) >> 8) & ~255) | ((56304) & 255)) } else {(56304)}))), 
instr_type: ((4) | ((0) << 13) | (if (((56304) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fucomip, 
opcode: (u64((if (((57320) & 65280) == 3840){ ((((57320) >> 8) & ~255) | ((57320) & 255)) } else {(57320)}))), 
instr_type: ((4) | ((0) << 13) | (if (((57320) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_fcomip, 
opcode: (u64((if (((57328) & 65280) == 3840){ ((((57328) >> 8) & ~255) | ((57328) & 255)) } else {(57328)}))), 
instr_type: ((4) | ((0) << 13) | (if (((57328) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_st, opt_st0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movd, 
opcode: (u64((if (((3950) & 65280) == 3840){ ((((3950) >> 8) & ~255) | ((3950) & 255)) } else {(3950)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3950) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg32, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movd, 
opcode: (u64((if (((3950) & 65280) == 3840){ ((((3950) >> 8) & ~255) | ((3950) & 255)) } else {(3950)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3950) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg64, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((3950) & 65280) == 3840){ ((((3950) >> 8) & ~255) | ((3950) & 255)) } else {(3950)}))), 
instr_type: ((8 | 512) | ((0) << 13) | (if (((3950) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_reg64, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((3951) & 65280) == 3840){ ((((3951) >> 8) & ~255) | ((3951) & 255)) } else {(3951)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3951) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmx, opt_mmx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movd, 
opcode: (u64((if (((3966) & 65280) == 3840){ ((((3966) >> 8) & ~255) | ((3966) & 255)) } else {(3966)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3966) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_mmxsse, opt_ea | opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movd, 
opcode: (u64((if (((3966) & 65280) == 3840){ ((((3966) >> 8) & ~255) | ((3966) & 255)) } else {(3966)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3966) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_mmxsse, opt_ea | opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((3967) & 65280) == 3840){ ((((3967) >> 8) & ~255) | ((3967) & 255)) } else {(3967)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3967) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_mmx, opt_ea | opt_mmx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((6688726) & 65280) == 3840){ ((((6688726) >> 8) & ~255) | ((6688726) & 255)) } else {(6688726)}))), 
instr_type: ((8) | ((0) << 13) | (if (((6688726) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_sse, opt_ea | opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((15929214) & 65280) == 3840){ ((((15929214) >> 8) & ~255) | ((15929214) & 255)) } else {(15929214)}))), 
instr_type: ((8) | ((0) << 13) | (if (((15929214) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movq, 
opcode: (u64((if (((3966) & 65280) == 3840){ ((((3966) >> 8) & ~255) | ((3966) & 255)) } else {(3966)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3966) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_mmxsse, opt_ea | opt_reg64]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_packssdw, 
opcode: (u64((if (((3947) & 65280) == 3840){ ((((3947) >> 8) & ~255) | ((3947) & 255)) } else {(3947)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3947) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_packsswb, 
opcode: (u64((if (((3939) & 65280) == 3840){ ((((3939) >> 8) & ~255) | ((3939) & 255)) } else {(3939)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3939) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_packuswb, 
opcode: (u64((if (((3943) & 65280) == 3840){ ((((3943) >> 8) & ~255) | ((3943) & 255)) } else {(3943)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3943) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddb, 
opcode: (u64((if (((4092) & 65280) == 3840){ ((((4092) >> 8) & ~255) | ((4092) & 255)) } else {(4092)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4092) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddw, 
opcode: (u64((if (((4093) & 65280) == 3840){ ((((4093) >> 8) & ~255) | ((4093) & 255)) } else {(4093)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4093) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddd, 
opcode: (u64((if (((4094) & 65280) == 3840){ ((((4094) >> 8) & ~255) | ((4094) & 255)) } else {(4094)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4094) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddsb, 
opcode: (u64((if (((4076) & 65280) == 3840){ ((((4076) >> 8) & ~255) | ((4076) & 255)) } else {(4076)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4076) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddsw, 
opcode: (u64((if (((4077) & 65280) == 3840){ ((((4077) >> 8) & ~255) | ((4077) & 255)) } else {(4077)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4077) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddusb, 
opcode: (u64((if (((4060) & 65280) == 3840){ ((((4060) >> 8) & ~255) | ((4060) & 255)) } else {(4060)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4060) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_paddusw, 
opcode: (u64((if (((4061) & 65280) == 3840){ ((((4061) >> 8) & ~255) | ((4061) & 255)) } else {(4061)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4061) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pand, 
opcode: (u64((if (((4059) & 65280) == 3840){ ((((4059) >> 8) & ~255) | ((4059) & 255)) } else {(4059)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4059) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pandn, 
opcode: (u64((if (((4063) & 65280) == 3840){ ((((4063) >> 8) & ~255) | ((4063) & 255)) } else {(4063)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4063) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpeqb, 
opcode: (u64((if (((3956) & 65280) == 3840){ ((((3956) >> 8) & ~255) | ((3956) & 255)) } else {(3956)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3956) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpeqw, 
opcode: (u64((if (((3957) & 65280) == 3840){ ((((3957) >> 8) & ~255) | ((3957) & 255)) } else {(3957)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3957) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpeqd, 
opcode: (u64((if (((3958) & 65280) == 3840){ ((((3958) >> 8) & ~255) | ((3958) & 255)) } else {(3958)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3958) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpgtb, 
opcode: (u64((if (((3940) & 65280) == 3840){ ((((3940) >> 8) & ~255) | ((3940) & 255)) } else {(3940)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3940) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpgtw, 
opcode: (u64((if (((3941) & 65280) == 3840){ ((((3941) >> 8) & ~255) | ((3941) & 255)) } else {(3941)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3941) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pcmpgtd, 
opcode: (u64((if (((3942) & 65280) == 3840){ ((((3942) >> 8) & ~255) | ((3942) & 255)) } else {(3942)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3942) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pmaddwd, 
opcode: (u64((if (((4085) & 65280) == 3840){ ((((4085) >> 8) & ~255) | ((4085) & 255)) } else {(4085)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4085) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pmulhw, 
opcode: (u64((if (((4069) & 65280) == 3840){ ((((4069) >> 8) & ~255) | ((4069) & 255)) } else {(4069)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4069) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pmullw, 
opcode: (u64((if (((4053) & 65280) == 3840){ ((((4053) >> 8) & ~255) | ((4053) & 255)) } else {(4053)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4053) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_por, 
opcode: (u64((if (((4075) & 65280) == 3840){ ((((4075) >> 8) & ~255) | ((4075) & 255)) } else {(4075)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4075) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psllw, 
opcode: (u64((if (((4081) & 65280) == 3840){ ((((4081) >> 8) & ~255) | ((4081) & 255)) } else {(4081)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4081) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psllw, 
opcode: (u64((if (((3953) & 65280) == 3840){ ((((3953) >> 8) & ~255) | ((3953) & 255)) } else {(3953)}))), 
instr_type: ((8) | ((6) << 13) | (if (((3953) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pslld, 
opcode: (u64((if (((4082) & 65280) == 3840){ ((((4082) >> 8) & ~255) | ((4082) & 255)) } else {(4082)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4082) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pslld, 
opcode: (u64((if (((3954) & 65280) == 3840){ ((((3954) >> 8) & ~255) | ((3954) & 255)) } else {(3954)}))), 
instr_type: ((8) | ((6) << 13) | (if (((3954) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psllq, 
opcode: (u64((if (((4083) & 65280) == 3840){ ((((4083) >> 8) & ~255) | ((4083) & 255)) } else {(4083)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4083) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psllq, 
opcode: (u64((if (((3955) & 65280) == 3840){ ((((3955) >> 8) & ~255) | ((3955) & 255)) } else {(3955)}))), 
instr_type: ((8) | ((6) << 13) | (if (((3955) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psraw, 
opcode: (u64((if (((4065) & 65280) == 3840){ ((((4065) >> 8) & ~255) | ((4065) & 255)) } else {(4065)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4065) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psraw, 
opcode: (u64((if (((3953) & 65280) == 3840){ ((((3953) >> 8) & ~255) | ((3953) & 255)) } else {(3953)}))), 
instr_type: ((8) | ((4) << 13) | (if (((3953) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrad, 
opcode: (u64((if (((4066) & 65280) == 3840){ ((((4066) >> 8) & ~255) | ((4066) & 255)) } else {(4066)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4066) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrad, 
opcode: (u64((if (((3954) & 65280) == 3840){ ((((3954) >> 8) & ~255) | ((3954) & 255)) } else {(3954)}))), 
instr_type: ((8) | ((4) << 13) | (if (((3954) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrlw, 
opcode: (u64((if (((4049) & 65280) == 3840){ ((((4049) >> 8) & ~255) | ((4049) & 255)) } else {(4049)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4049) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrlw, 
opcode: (u64((if (((3953) & 65280) == 3840){ ((((3953) >> 8) & ~255) | ((3953) & 255)) } else {(3953)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3953) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrld, 
opcode: (u64((if (((4050) & 65280) == 3840){ ((((4050) >> 8) & ~255) | ((4050) & 255)) } else {(4050)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4050) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrld, 
opcode: (u64((if (((3954) & 65280) == 3840){ ((((3954) >> 8) & ~255) | ((3954) & 255)) } else {(3954)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3954) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrlq, 
opcode: (u64((if (((4051) & 65280) == 3840){ ((((4051) >> 8) & ~255) | ((4051) & 255)) } else {(4051)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4051) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psrlq, 
opcode: (u64((if (((3955) & 65280) == 3840){ ((((3955) >> 8) & ~255) | ((3955) & 255)) } else {(3955)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3955) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_im8, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubb, 
opcode: (u64((if (((4088) & 65280) == 3840){ ((((4088) >> 8) & ~255) | ((4088) & 255)) } else {(4088)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4088) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubw, 
opcode: (u64((if (((4089) & 65280) == 3840){ ((((4089) >> 8) & ~255) | ((4089) & 255)) } else {(4089)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4089) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubd, 
opcode: (u64((if (((4090) & 65280) == 3840){ ((((4090) >> 8) & ~255) | ((4090) & 255)) } else {(4090)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4090) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubsb, 
opcode: (u64((if (((4072) & 65280) == 3840){ ((((4072) >> 8) & ~255) | ((4072) & 255)) } else {(4072)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4072) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubsw, 
opcode: (u64((if (((4073) & 65280) == 3840){ ((((4073) >> 8) & ~255) | ((4073) & 255)) } else {(4073)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4073) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubusb, 
opcode: (u64((if (((4056) & 65280) == 3840){ ((((4056) >> 8) & ~255) | ((4056) & 255)) } else {(4056)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4056) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_psubusw, 
opcode: (u64((if (((4057) & 65280) == 3840){ ((((4057) >> 8) & ~255) | ((4057) & 255)) } else {(4057)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4057) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpckhbw, 
opcode: (u64((if (((3944) & 65280) == 3840){ ((((3944) >> 8) & ~255) | ((3944) & 255)) } else {(3944)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3944) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpckhwd, 
opcode: (u64((if (((3945) & 65280) == 3840){ ((((3945) >> 8) & ~255) | ((3945) & 255)) } else {(3945)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3945) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpckhdq, 
opcode: (u64((if (((3946) & 65280) == 3840){ ((((3946) >> 8) & ~255) | ((3946) & 255)) } else {(3946)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3946) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpcklbw, 
opcode: (u64((if (((3936) & 65280) == 3840){ ((((3936) >> 8) & ~255) | ((3936) & 255)) } else {(3936)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3936) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpcklwd, 
opcode: (u64((if (((3937) & 65280) == 3840){ ((((3937) >> 8) & ~255) | ((3937) & 255)) } else {(3937)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3937) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_punpckldq, 
opcode: (u64((if (((3938) & 65280) == 3840){ ((((3938) >> 8) & ~255) | ((3938) & 255)) } else {(3938)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3938) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pxor, 
opcode: (u64((if (((4079) & 65280) == 3840){ ((((4079) >> 8) & ~255) | ((4079) & 255)) } else {(4079)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4079) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movups, 
opcode: (u64((if (((3856) & 65280) == 3840){ ((((3856) >> 8) & ~255) | ((3856) & 255)) } else {(3856)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3856) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg32, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movups, 
opcode: (u64((if (((3857) & 65280) == 3840){ ((((3857) >> 8) & ~255) | ((3857) & 255)) } else {(3857)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3857) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_sse, opt_ea | opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movaps, 
opcode: (u64((if (((3880) & 65280) == 3840){ ((((3880) >> 8) & ~255) | ((3880) & 255)) } else {(3880)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3880) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg32, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movaps, 
opcode: (u64((if (((3881) & 65280) == 3840){ ((((3881) >> 8) & ~255) | ((3881) & 255)) } else {(3881)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3881) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_sse, opt_ea | opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movhps, 
opcode: (u64((if (((3862) & 65280) == 3840){ ((((3862) >> 8) & ~255) | ((3862) & 255)) } else {(3862)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3862) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_reg32, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_movhps, 
opcode: (u64((if (((3863) & 65280) == 3840){ ((((3863) >> 8) & ~255) | ((3863) & 255)) } else {(3863)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3863) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_sse, opt_ea | opt_reg32]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_addps, 
opcode: (u64((if (((3928) & 65280) == 3840){ ((((3928) >> 8) & ~255) | ((3928) & 255)) } else {(3928)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3928) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cvtpi2ps, 
opcode: (u64((if (((3882) & 65280) == 3840){ ((((3882) >> 8) & ~255) | ((3882) & 255)) } else {(3882)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3882) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmx, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cvtps2pi, 
opcode: (u64((if (((3885) & 65280) == 3840){ ((((3885) >> 8) & ~255) | ((3885) & 255)) } else {(3885)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3885) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_mmx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_cvttps2pi, 
opcode: (u64((if (((3884) & 65280) == 3840){ ((((3884) >> 8) & ~255) | ((3884) & 255)) } else {(3884)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3884) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_mmx]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_divps, 
opcode: (u64((if (((3934) & 65280) == 3840){ ((((3934) >> 8) & ~255) | ((3934) & 255)) } else {(3934)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3934) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_maxps, 
opcode: (u64((if (((3935) & 65280) == 3840){ ((((3935) >> 8) & ~255) | ((3935) & 255)) } else {(3935)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3935) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_minps, 
opcode: (u64((if (((3933) & 65280) == 3840){ ((((3933) >> 8) & ~255) | ((3933) & 255)) } else {(3933)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3933) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_mulps, 
opcode: (u64((if (((3929) & 65280) == 3840){ ((((3929) >> 8) & ~255) | ((3929) & 255)) } else {(3929)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3929) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pavgb, 
opcode: (u64((if (((4064) & 65280) == 3840){ ((((4064) >> 8) & ~255) | ((4064) & 255)) } else {(4064)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4064) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pavgw, 
opcode: (u64((if (((4067) & 65280) == 3840){ ((((4067) >> 8) & ~255) | ((4067) & 255)) } else {(4067)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4067) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pmaxsw, 
opcode: (u64((if (((4078) & 65280) == 3840){ ((((4078) >> 8) & ~255) | ((4078) & 255)) } else {(4078)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4078) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pmaxub, 
opcode: (u64((if (((4062) & 65280) == 3840){ ((((4062) >> 8) & ~255) | ((4062) & 255)) } else {(4062)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4062) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pminsw, 
opcode: (u64((if (((4074) & 65280) == 3840){ ((((4074) >> 8) & ~255) | ((4074) & 255)) } else {(4074)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4074) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_pminub, 
opcode: (u64((if (((4058) & 65280) == 3840){ ((((4058) >> 8) & ~255) | ((4058) & 255)) } else {(4058)}))), 
instr_type: ((8) | ((0) << 13) | (if (((4058) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_mmxsse, opt_mmxsse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_rcpss, 
opcode: (u64((if (((3923) & 65280) == 3840){ ((((3923) >> 8) & ~255) | ((3923) & 255)) } else {(3923)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3923) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_rsqrtps, 
opcode: (u64((if (((3922) & 65280) == 3840){ ((((3922) >> 8) & ~255) | ((3922) & 255)) } else {(3922)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3922) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sqrtps, 
opcode: (u64((if (((3921) & 65280) == 3840){ ((((3921) >> 8) & ~255) | ((3921) & 255)) } else {(3921)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3921) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_subps, 
opcode: (u64((if (((3932) & 65280) == 3840){ ((((3932) >> 8) & ~255) | ((3932) & 255)) } else {(3932)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3932) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 2, 
op_type: [opt_ea | opt_sse, opt_sse]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_prefetchnta, 
opcode: (u64((if (((3864) & 65280) == 3840){ ((((3864) >> 8) & ~255) | ((3864) & 255)) } else {(3864)}))), 
instr_type: ((8) | ((0) << 13) | (if (((3864) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_prefetcht0, 
opcode: (u64((if (((3864) & 65280) == 3840){ ((((3864) >> 8) & ~255) | ((3864) & 255)) } else {(3864)}))), 
instr_type: ((8) | ((1) << 13) | (if (((3864) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_prefetcht1, 
opcode: (u64((if (((3864) & 65280) == 3840){ ((((3864) >> 8) & ~255) | ((3864) & 255)) } else {(3864)}))), 
instr_type: ((8) | ((2) << 13) | (if (((3864) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_prefetcht2, 
opcode: (u64((if (((3864) & 65280) == 3840){ ((((3864) >> 8) & ~255) | ((3864) & 255)) } else {(3864)}))), 
instr_type: ((8) | ((3) << 13) | (if (((3864) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_prefetchw, 
opcode: (u64((if (((3853) & 65280) == 3840){ ((((3853) >> 8) & ~255) | ((3853) & 255)) } else {(3853)}))), 
instr_type: ((8) | ((1) << 13) | (if (((3853) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_lfence, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((5) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_mfence, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((6) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_sfence, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((7) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 0, 
op_type: [0]!

}
, ASMInstr {
sym: Tcc_token.tok_asm_clflush, 
opcode: (u64((if (((4014) & 65280) == 3840){ ((((4014) >> 8) & ~255) | ((4014) & 255)) } else {(4014)}))), 
instr_type: ((8) | ((7) << 13) | (if (((4014) & 65280) == 3840){ 256 } else {0})), 
nb_ops: 1, 
op_type: [opt_ea]!

}
, ASMInstr {
sym: 0, 
}
]!

)

[export:'op0_codes']
const (
op0_codes   = [248, 252, 250, 3846, 245, 159, 158, 156, 157, 156, 157, 249, 253, 251, 55, 63, 39, 47, 54538, 54282, 26264, 26265, 152, 153, 26264, 152, 26265, 153, 18585, 204, 206, 207, 4010, 244, 155, 144, 62352, 215, 240, 243, 243, 243, 242, 242, 3848, 3849, 4002, 3888, 3889, 3890, 3891, 3845, 3847, 3851, 201, 195, 195, 203, 56041, 55780, 55781, 55784, 55785, 55786, 55787, 55788, 55789, 55790, 55792, 55793, 55794, 55795, 55796, 55797, 55798, 55799, 55800, 55801, 55802, 55803, 55804, 55805, 55806, 55807, 55776, 55777, 56291, 56290, 55760, 155, 55753, 57312, 3959]!

)

fn tcc_basename(name &i8) &i8 {
	p := C.strchr(name, 0)
	for p > name && !(p [-1]  == `/`) {
	p --$
	}
	return p
}

fn tcc_fileextension(name &i8) &i8 {
	b := tcc_basename(name)
	e := C.strrchr(b, `.`)
	return if e{ e } else {C.strchr(b, 0)}
}

fn tcc_strdup(str &i8) &i8 {
	ptr := &i8(0)
	ptr = tcc_malloc(C.strlen(str) + 1)
	strcpy(ptr, str)
	return ptr
}

@[c2v_variadic]
fn tcc_error(fmt &i8)  {
	s1 := tcc_state
	ap := Va_list{}
	__builtin_va_start(ap, fmt)
	error1(s1, 0, fmt, ap)
	__builtin_va_end(ap)
	if s1.error_set_jmp_enabled {
		longjmp(s1.error_jmp_buf, 1)
	}
	else {
		C.exit(1)
	}
}

fn tcc_new() &TCCState {
	s := &TCCState(0)
	tcc_cleanup()
	s = tcc_mallocz(sizeof(TCCState))
	if !s {
	return (voidptr(0))
	}
	tcc_state = s
	nb_states ++$
	s.nocommon = 1
	s.dollars_in_identifiers = 1
	s.cversion = 199901
	s.warn_implicit_function_declaration = 1
	s.ms_extensions = 1
	tcc_set_lib_path(s, c'/usr/local/lib/tcc')
	tccelf_new(s)
	tccpp_new(s)
	define_push(Tcc_token.tok___line__, 0, (voidptr(0)), (voidptr(0)))
	define_push(Tcc_token.tok___file__, 0, (voidptr(0)), (voidptr(0)))
	define_push(Tcc_token.tok___date__, 0, (voidptr(0)), (voidptr(0)))
	define_push(Tcc_token.tok___time__, 0, (voidptr(0)), (voidptr(0)))
	define_push(Tcc_token.tok___counter__, 0, (voidptr(0)), (voidptr(0)))
	{
		buffer := [32]i8{}
		a := 0
		b := 0
		c := 0
		
		C.sscanf(c'0.9.27', c'%d.%d.%d', &a, &b, &c)
		sprintf(buffer, c'%d', a * 10000 + b * 100 + c)
		tcc_define_symbol(s, c'__TINYC__', buffer)
	}
	tcc_define_symbol(s, c'__STDC__', (voidptr(0)))
	tcc_define_symbol(s, c'__STDC_VERSION__', c'199901L')
	tcc_define_symbol(s, c'__STDC_HOSTED__', (voidptr(0)))
	tcc_define_symbol(s, c'__x86_64__', (voidptr(0)))
	tcc_define_symbol(s, c'__unix__', (voidptr(0)))
	tcc_define_symbol(s, c'__unix', (voidptr(0)))
	tcc_define_symbol(s, c'unix', (voidptr(0)))
	tcc_define_symbol(s, c'__linux__', (voidptr(0)))
	tcc_define_symbol(s, c'__linux', (voidptr(0)))
	tcc_define_symbol(s, c'__SIZE_TYPE__', c'unsigned long')
	tcc_define_symbol(s, c'__PTRDIFF_TYPE__', c'long')
	tcc_define_symbol(s, c'__LP64__', (voidptr(0)))
	tcc_define_symbol(s, c'__SIZEOF_POINTER__', if 8 == 4{ c'4' } else {c'8'})
	tcc_define_symbol(s, c'__WCHAR_TYPE__', c'int')
	tcc_define_symbol(s, c'__WINT_TYPE__', c'unsigned int')
	tcc_define_symbol(s, c'__REDIRECT(name, proto, alias)', c'name proto __asm__ (#alias)')
	tcc_define_symbol(s, c'__REDIRECT_NTH(name, proto, alias)', c'name proto __asm__ (#alias) __THROW')
	tcc_define_symbol(s, c'__builtin_extract_return_addr(x)', c'x')
	return s
}

fn tcc_delete(s1 &TCCState)  {
	tcc_cleanup()
	tccelf_delete(s1)
	dynarray_reset(&s1.library_paths, &s1.nb_library_paths)
	dynarray_reset(&s1.crt_paths, &s1.nb_crt_paths)
	dynarray_reset(&s1.cached_includes, &s1.nb_cached_includes)
	dynarray_reset(&s1.include_paths, &s1.nb_include_paths)
	dynarray_reset(&s1.sysinclude_paths, &s1.nb_sysinclude_paths)
	dynarray_reset(&s1.cmd_include_files, &s1.nb_cmd_include_files)
	tcc_free(s1.tcc_lib_path)
	tcc_free(s1.soname)
	tcc_free(s1.rpath)
	tcc_free(s1.init_symbol)
	tcc_free(s1.fini_symbol)
	tcc_free(s1.outfile)
	tcc_free(s1.deps_outfile)
	dynarray_reset(&s1.files, &s1.nb_files)
	dynarray_reset(&s1.target_deps, &s1.nb_target_deps)
	dynarray_reset(&s1.pragma_libs, &s1.nb_pragma_libs)
	dynarray_reset(&s1.argv, &s1.argc)
	tcc_run_free(s1)
	tcc_free(s1)
	if 0 == nb_states --$ {
	tcc_memcheck()
	}
}

fn tcc_set_output_type(s &TCCState, output_type int) int {
	s.output_type = output_type
	if output_type == 4 {
	s.output_format = 0
	}
	if s.char_is_unsigned {
	tcc_define_symbol(s, c'__CHAR_UNSIGNED__', (voidptr(0)))
	}
	if !s.nostdinc {
		tcc_add_sysinclude_path(s, c'{B}/include:/usr/local/include:/usr/include')
	}
	if s.do_bounds_check {
		tccelf_bounds_new(s)
		tcc_define_symbol(s, c'__BOUNDS_CHECKING_ON', (voidptr(0)))
	}
	if s.do_debug {
		tccelf_stab_new(s)
	}
	tcc_add_library_path(s, c'/usr/lib:/lib:/usr/local/lib')
	tcc_split_path(s, &s.crt_paths, &s.nb_crt_paths, c'/usr/lib')
	if (output_type == 2 || output_type == 3) && !s.nostdlib {
		if output_type != 3 {
		tcc_add_crt(s, c'crt1.o')
		}
		tcc_add_crt(s, c'crti.o')
	}
	return 0
}

fn tcc_add_include_path(s &TCCState, pathname &i8) int {
	tcc_split_path(s, &s.include_paths, &s.nb_include_paths, pathname)
	return 0
}

fn tcc_add_sysinclude_path(s &TCCState, pathname &i8) int {
	tcc_split_path(s, &s.sysinclude_paths, &s.nb_sysinclude_paths, pathname)
	return 0
}

fn tcc_add_file(s &TCCState, filename &i8) int {
	filetype := s.filetype
	if 0 == (filetype & (15 | 64)) {
		ext := tcc_fileextension(filename)
		if ext [0]  {
			ext ++
			if !C.strcmp(ext, c'S') {
			filetype = 4
			}
			else if !C.strcmp(ext, c's') {
			filetype = 2
			}
			else if !C.strcmp(ext, c'c') || !C.strcmp(ext, c'i') {
			filetype = 1
			}
			else { // 3
			filetype |= 64
}
		}
		else {
			filetype = 1
		}
	}
	return tcc_add_file_internal(s, filename, filetype | 16)
}

fn tcc_add_library_path(s &TCCState, pathname &i8) int {
	tcc_split_path(s, &s.library_paths, &s.nb_library_paths, pathname)
	return 0
}

fn tcc_add_library(s &TCCState, libraryname &i8) int {
	libs := [c'%s/lib%s.so', c'%s/lib%s.a', (voidptr(0))]!
	
	pp := if s.static_link{ libs + 1 } else {libs}
	flags := s.filetype & 128
	for *pp {
		if 0 == tcc_add_library_internal(s, *pp, libraryname, flags, s.library_paths, s.nb_library_paths) {
		return 0
		}
		pp ++$
	}
	return -1
}

fn tcc_add_library_err(s &TCCState, libname &i8) int {
	ret := tcc_add_library(s, libname)
	if ret < 0 {
	tcc_error_noabort(c"library '%s' not found", libname)
	}
	return ret
}

struct FlagDef { 
	offset u16
	flags u16
	name &i8
}
struct TCCOption { 
	name &i8
	index u16
	flags u16
}

const ( // empty enum
	tcc_option_help = 0
	tcc_option_help2 = 1
	tcc_option_v = 2
	tcc_option_i = 3
	tcc_option_d = 4
	tcc_option_u = 5
	tcc_option_p = 6
	tcc_option_l = 7
	tcc_option_b = 8

	tcc_option_bench = 10
	tcc_option_bt = 11

	tcc_option_g = 13
	tcc_option_c = 14
	tcc_option_dumpversion = 15

	tcc_option_static = 17
	tcc_option_std = 18
	tcc_option_shared = 19
	tcc_option_soname = 20
	tcc_option_o = 21
	tcc_option_r = 22
	tcc_option_s = 23
	tcc_option_traditional = 24
	tcc_option_wl = 25
	tcc_option_wp = 26
	tcc_option_w = 27

	tcc_option_mfloat_abi = 29
	tcc_option_m = 30
	tcc_option_f = 31
	tcc_option_isystem = 32
	tcc_option_iwithprefix = 33
	tcc_option_include = 34
	tcc_option_nostdinc = 35
	tcc_option_nostdlib = 36
	tcc_option_print_search_dirs = 37
	tcc_option_rdynamic = 38
	tcc_option_param = 39
	tcc_option_pedantic = 40
	tcc_option_pthread = 41
	tcc_option_run = 42

	tcc_option_pipe = 44
	tcc_option_e = 45
	tcc_option_md = 46
	tcc_option_mf = 47
	tcc_option_x = 48
	tcc_option_ar = 49
	tcc_option_impdef = 50
)

[export:'tcc_options']
const (
tcc_options   = [TCCOption {
name: c'h', 
index: tcc_option_help, 
flags: 0
}
, TCCOption {
name: c'-help', 
index: tcc_option_help, 
flags: 0
}
, TCCOption {
name: c'?', 
index: tcc_option_help, 
flags: 0
}
, TCCOption {
name: c'hh', 
index: tcc_option_help2, 
flags: 0
}
, TCCOption {
name: c'v', 
index: tcc_option_v, 
flags: 1 | 2
}
, TCCOption {
name: c'I', 
index: tcc_option_i, 
flags: 1
}
, TCCOption {
name: c'D', 
index: tcc_option_d, 
flags: 1
}
, TCCOption {
name: c'U', 
index: tcc_option_u, 
flags: 1
}
, TCCOption {
name: c'P', 
index: tcc_option_p, 
flags: 1 | 2
}
, TCCOption {
name: c'L', 
index: tcc_option_l, 
flags: 1
}
, TCCOption {
name: c'B', 
index: tcc_option_b, 
flags: 1
}
, TCCOption {
name: c'l', 
index: tcc_option_l, 
flags: 1
}
, TCCOption {
name: c'bench', 
index: tcc_option_bench, 
flags: 0
}
, TCCOption {
name: c'bt', 
index: tcc_option_bt, 
flags: 1
}
, TCCOption {
name: c'b', 
index: tcc_option_b, 
flags: 0
}
, TCCOption {
name: c'g', 
index: tcc_option_g, 
flags: 1 | 2
}
, TCCOption {
name: c'c', 
index: tcc_option_c, 
flags: 0
}
, TCCOption {
name: c'dumpversion', 
index: tcc_option_dumpversion, 
flags: 0
}
, TCCOption {
name: c'd', 
index: tcc_option_d, 
flags: 1 | 2
}
, TCCOption {
name: c'static', 
index: tcc_option_static, 
flags: 0
}
, TCCOption {
name: c'std', 
index: tcc_option_std, 
flags: 1 | 2
}
, TCCOption {
name: c'shared', 
index: tcc_option_shared, 
flags: 0
}
, TCCOption {
name: c'soname', 
index: tcc_option_soname, 
flags: 1
}
, TCCOption {
name: c'o', 
index: tcc_option_o, 
flags: 1
}
, TCCOption {
name: c'-param', 
index: tcc_option_param, 
flags: 1
}
, TCCOption {
name: c'pedantic', 
index: tcc_option_pedantic, 
flags: 0
}
, TCCOption {
name: c'pthread', 
index: tcc_option_pthread, 
flags: 0
}
, TCCOption {
name: c'run', 
index: tcc_option_run, 
flags: 1 | 2
}
, TCCOption {
name: c'rdynamic', 
index: tcc_option_rdynamic, 
flags: 0
}
, TCCOption {
name: c'r', 
index: tcc_option_r, 
flags: 0
}
, TCCOption {
name: c's', 
index: tcc_option_s, 
flags: 0
}
, TCCOption {
name: c'traditional', 
index: tcc_option_traditional, 
flags: 0
}
, TCCOption {
name: c'Wl,', 
index: tcc_option_wl, 
flags: 1 | 2
}
, TCCOption {
name: c'Wp,', 
index: tcc_option_wp, 
flags: 1 | 2
}
, TCCOption {
name: c'W', 
index: tcc_option_w, 
flags: 1 | 2
}
, TCCOption {
name: c'O', 
index: tcc_option_o, 
flags: 1 | 2
}
, TCCOption {
name: c'm', 
index: tcc_option_m, 
flags: 1 | 2
}
, TCCOption {
name: c'f', 
index: tcc_option_f, 
flags: 1 | 2
}
, TCCOption {
name: c'isystem', 
index: tcc_option_isystem, 
flags: 1
}
, TCCOption {
name: c'include', 
index: tcc_option_include, 
flags: 1
}
, TCCOption {
name: c'nostdinc', 
index: tcc_option_nostdinc, 
flags: 0
}
, TCCOption {
name: c'nostdlib', 
index: tcc_option_nostdlib, 
flags: 0
}
, TCCOption {
name: c'print-search-dirs', 
index: tcc_option_print_search_dirs, 
flags: 0
}
, TCCOption {
name: c'w', 
index: tcc_option_w, 
flags: 0
}
, TCCOption {
name: c'pipe', 
index: tcc_option_pipe, 
flags: 0
}
, TCCOption {
name: c'E', 
index: tcc_option_e, 
flags: 0
}
, TCCOption {
name: c'MD', 
index: tcc_option_md, 
flags: 0
}
, TCCOption {
name: c'MF', 
index: tcc_option_mf, 
flags: 1
}
, TCCOption {
name: c'x', 
index: tcc_option_x, 
flags: 1
}
, TCCOption {
name: c'ar', 
index: tcc_option_ar, 
flags: 0
}
, TCCOption {
name: (voidptr(0)), 
index: 0, 
flags: 0
}
]!

)

[export:'options_W']
const (
options_W   = [FlagDef {
offset: 0, 
flags: 0, 
name: c'all'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).warn_unsupported)), 
flags: 0, 
name: c'unsupported'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).warn_write_strings)), 
flags: 0, 
name: c'write-strings'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).warn_error)), 
flags: 0, 
name: c'error'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).warn_gcc_compat)), 
flags: 0, 
name: c'gcc-compat'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).warn_implicit_function_declaration)), 
flags: 1, 
name: c'implicit-function-declaration'
}
, FlagDef {
offset: 0, 
flags: 0, 
name: (voidptr(0))
}
]!

)

[export:'options_f']
const (
options_f   = [FlagDef {
offset: (usize(&(&TCCState(0)).char_is_unsigned)), 
flags: 0, 
name: c'unsigned-char'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).char_is_unsigned)), 
flags: 2, 
name: c'signed-char'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).nocommon)), 
flags: 2, 
name: c'common'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).leading_underscore)), 
flags: 0, 
name: c'leading-underscore'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).ms_extensions)), 
flags: 0, 
name: c'ms-extensions'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).dollars_in_identifiers)), 
flags: 0, 
name: c'dollars-in-identifiers'
}
, FlagDef {
offset: 0, 
flags: 0, 
name: (voidptr(0))
}
]!

)

[export:'options_m']
const (
options_m   = [FlagDef {
offset: (usize(&(&TCCState(0)).ms_bitfields)), 
flags: 0, 
name: c'ms-bitfields'
}
, FlagDef {
offset: (usize(&(&TCCState(0)).nosse)), 
flags: 2, 
name: c'sse'
}
, FlagDef {
offset: 0, 
flags: 0, 
name: (voidptr(0))
}
]!

)

fn tcc_parse_args(s &TCCState, pargc &int, pargv &&&i8, optind int) int {
	popt := &TCCOption(0)
	optarg := &i8(0)
	r := &i8(0)
	
	run := (voidptr(0))
	last_o := -1
	x := 0
	linker_arg := CString{}
	tool := 0
arg_start := 0
noaction := optind

	argv := *pargv
	argc := *pargc
	cstr_new(&linker_arg)
	for optind < argc {
		r = argv [optind] 
		if r [0]  == `@` && r [1]  != ` ` {
			args_parser_listfile(s, r + 1, optind, &argc, &argv)
			continue
			
		}
		optind ++
		if tool {
			if r [0]  == `-` && r [1]  == `v` && r [2]  == 0 {
			s.verbose ++$
			}
			continue
			
		}
		// RRRREG reparse id=0x7fffc1f88b48
		reparse: 
		if r [0]  != `-` || r [1]  == ` ` {
			if r [0]  != `@` {
			args_parser_add_file(s, r, s.filetype)
			}
			if run {
				tcc_set_options(s, run)
				arg_start = optind - 1
				break
				
			}
			continue
			
		}
		for popt = tcc_options ;  ; popt ++ {
			p1 := popt.name
			r1 := r + 1
			if p1 == (voidptr(0)) {
			tcc_error(c"invalid option -- '%s'", r)
			}
			if !strstart(p1, &r1) {
			continue
			
			}
			optarg = r1
			if popt.flags & 1 {
				if *r1 == ` ` && !(popt.flags & 2) {
					if optind >= argc {
					// RRRREG arg_err id=0x7fffc1f89688
					arg_err: 
					tcc_error(c"argument to '%s' is missing", r)
					}
					optarg = argv [optind ++] 
				}
			}
			else if *r1 != ` ` {
			continue
			
			}
			break
			
		}
		match (popt.index) {
		 tcc_option_help{ // case comp body kind=ReturnStmt is_enum=true
		return 1
		}
		 tcc_option_help2{ // case comp body kind=ReturnStmt is_enum=true
		return 2
		}
		 tcc_option_i{ // case comp body kind=CallExpr is_enum=true
		tcc_add_include_path(s, optarg)
		
		}
		 tcc_option_d{ // case comp body kind=CallExpr is_enum=true
		parse_option_d(s, optarg)
		
		}
		 tcc_option_u{ // case comp body kind=CallExpr is_enum=true
		tcc_undefine_symbol(s, optarg)
		
		}
		 tcc_option_l{ // case comp body kind=CallExpr is_enum=true
		tcc_add_library_path(s, optarg)
		
		}
		 tcc_option_b{ // case comp body kind=CallExpr is_enum=true
		tcc_set_lib_path(s, optarg)
		
		}
		 tcc_option_l{ // case comp body kind=CallExpr is_enum=true
		args_parser_add_file(s, optarg, 8 | (s.filetype & ~(15 | 64)))
		s.nb_libraries ++
		
		}
		 tcc_option_pthread{ // case comp body kind=CallExpr is_enum=true
		parse_option_d(s, c'_REENTRANT')
		s.option_pthread = 1
		
		}
		 tcc_option_bench{ // case comp body kind=BinaryOperator is_enum=true
		s.do_bench = 1
		
		}
		 tcc_option_bt{ // case comp body kind=CallExpr is_enum=true
		tcc_set_num_callers(C.atoi(optarg))
		
		}
		 tcc_option_b{ // case comp body kind=BinaryOperator is_enum=true
		s.do_bounds_check = 1
		s.do_debug = 1
		
		}
		 tcc_option_g{ // case comp body kind=BinaryOperator is_enum=true
		s.do_debug = 1
		
		}
		 tcc_option_c{ // case comp body kind=BinaryOperator is_enum=true
		x = 4
		// RRRREG set_output_type id=0x7fffc1f8afb0
		set_output_type: 
		if s.output_type {
		tcc_warning(c'-%s: overriding compiler action already specified', popt.name)
		}
		s.output_type = x
		
		}
		 tcc_option_d{ // case comp body kind=IfStmt is_enum=true
		if *optarg == `D` {
		s.dflag = 3
		}
		else if *optarg == `M` {
		s.dflag = 7
		}
		else if *optarg == `t` {
		s.dflag = 16
		}
		else if isnum(*optarg) {
		g_debug = C.atoi(optarg)
		}
		else { // 3
		goto unsupported_option // id: 0x7fffc1f8b768
		
}
		
		}
		 tcc_option_static{ // case comp body kind=BinaryOperator is_enum=true
		s.static_link = 1
		
		}
		 tcc_option_std{ // case comp body kind=IfStmt is_enum=true
		if *optarg == `=` {
			if C.strcmp(optarg, c'=c11') == 0 {
				tcc_undefine_symbol(s, c'__STDC_VERSION__')
				tcc_define_symbol(s, c'__STDC_VERSION__', c'201112L')
				tcc_define_symbol(s, c'__STDC_NO_ATOMICS__', c'1')
				tcc_define_symbol(s, c'__STDC_NO_COMPLEX__', c'1')
				tcc_define_symbol(s, c'__STDC_NO_THREADS__', c'1')
				tcc_define_symbol(s, c'__STDC_UTF_16__', c'1')
				tcc_define_symbol(s, c'__STDC_UTF_32__', c'1')
				s.cversion = 201112
			}
		}
		
		}
		 tcc_option_shared{ // case comp body kind=BinaryOperator is_enum=true
		x = 3
		goto set_output_type // id: 0x7fffc1f8afb0
		}
		 tcc_option_soname{ // case comp body kind=BinaryOperator is_enum=true
		s.soname = tcc_strdup(optarg)
		
		}
		 tcc_option_o{ // case comp body kind=IfStmt is_enum=true
		if s.outfile {
			tcc_warning(c'multiple -o option')
			tcc_free(s.outfile)
		}
		s.outfile = tcc_strdup(optarg)
		
		}
		 tcc_option_r{ // case comp body kind=BinaryOperator is_enum=true
		s.option_r = 1
		x = 4
		goto set_output_type // id: 0x7fffc1f8afb0
		}
		 tcc_option_isystem{ // case comp body kind=CallExpr is_enum=true
		tcc_add_sysinclude_path(s, optarg)
		
		}
		 tcc_option_include{ // case comp body kind=CallExpr is_enum=true
		dynarray_add(&s.cmd_include_files, &s.nb_cmd_include_files, tcc_strdup(optarg))
		
		}
		 tcc_option_nostdinc{ // case comp body kind=BinaryOperator is_enum=true
		s.nostdinc = 1
		
		}
		 tcc_option_nostdlib{ // case comp body kind=BinaryOperator is_enum=true
		s.nostdlib = 1
		
		}
		 tcc_option_run{ // case comp body kind=BinaryOperator is_enum=true
		run = optarg
		x = 1
		goto set_output_type // id: 0x7fffc1f8afb0
		}
		 tcc_option_v{ // case comp body kind=DoStmt is_enum=true
		for {
		s.verbose
		// while()
		if ! (*optarg ++ == `v` ) { break }
		}
		noaction ++$
		
		}
		 tcc_option_f{ // case comp body kind=IfStmt is_enum=true
		if set_flag(s, options_f, optarg) < 0 {
		goto unsupported_option // id: 0x7fffc1f8b768
		}
		
		}
		 tcc_option_m{ // case comp body kind=IfStmt is_enum=true
		if set_flag(s, options_m, optarg) < 0 {
			if x = C.atoi(optarg) , x != 32 && x != 64 {
			goto unsupported_option // id: 0x7fffc1f8b768
			}
			if 8 != x / 8 {
			return x
			}
			noaction ++$
		}
		
		}
		 tcc_option_w{ // case comp body kind=IfStmt is_enum=true
		if set_flag(s, options_W, optarg) < 0 {
		goto unsupported_option // id: 0x7fffc1f8b768
		}
		
		}
		 tcc_option_w{ // case comp body kind=BinaryOperator is_enum=true
		s.warn_none = 1
		
		}
		 tcc_option_rdynamic{ // case comp body kind=BinaryOperator is_enum=true
		s.rdynamic = 1
		
		}
		 tcc_option_wl{ // case comp body kind=IfStmt is_enum=true
		if linker_arg.size {
		linker_arg.size --$ , cstr_ccat(&linker_arg, `,`)
		}
		cstr_cat(&linker_arg, optarg, 0)
		if tcc_set_linker(s, linker_arg.data) {
		cstr_free(&linker_arg)
		}
		
		}
		 tcc_option_wp{ // case comp body kind=BinaryOperator is_enum=true
		r = optarg
		goto reparse // id: 0x7fffc1f88b48
		}
		 tcc_option_e{ // case comp body kind=BinaryOperator is_enum=true
		x = 5
		goto set_output_type // id: 0x7fffc1f8afb0
		}
		 tcc_option_p{ // case comp body kind=BinaryOperator is_enum=true
		s.Pflag = C.atoi(optarg) + 1
		
		}
		 tcc_option_md{ // case comp body kind=BinaryOperator is_enum=true
		s.gen_deps = 1
		
		}
		 tcc_option_mf{ // case comp body kind=BinaryOperator is_enum=true
		s.deps_outfile = tcc_strdup(optarg)
		
		}
		 tcc_option_dumpversion{ // case comp body kind=CallExpr is_enum=true
		C.printf(c'%s\n', c'0.9.27')
		C.exit(0)
		
		}
		 tcc_option_x{ // case comp body kind=BinaryOperator is_enum=true
		x = 0
		if *optarg == `c` {
		x = 1
		}
		else if *optarg == `a` {
		x = 4
		}
		else if *optarg == `b` {
		x = 64
		}
		else if *optarg == `n` {
		x = 0
		}
		else { // 3
		tcc_warning(c"unsupported language '%s'", optarg)
}
		s.filetype = x | (s.filetype & ~(15 | 64))
		
		}
		 tcc_option_o{ // case comp body kind=BinaryOperator is_enum=true
		last_o = C.atoi(optarg)
		
		}
		 tcc_option_print_search_dirs{ // case comp body kind=BinaryOperator is_enum=true
		x = 4
		goto extra_action // id: 0x7fffc1f8fbf8
		}
		 tcc_option_impdef{ // case comp body kind=BinaryOperator is_enum=true
		x = 6
		goto extra_action // id: 0x7fffc1f8fbf8
		}
		 tcc_option_ar{ // case comp body kind=BinaryOperator is_enum=true
		x = 5
		// RRRREG extra_action id=0x7fffc1f8fbf8
		extra_action: 
		arg_start = optind - 1
		if arg_start != noaction {
		tcc_error(c'cannot parse %s here', r)
		}
		tool = x
		
		}
		 tcc_option_traditional, tcc_option_pedantic, tcc_option_pipe, tcc_option_s{
		
		
		}
		else {
		// RRRREG unsupported_option id=0x7fffc1f8b768
		unsupported_option: 
		if s.warn_unsupported {
		tcc_warning(c"unsupported option '%s'", r)
		}
		}
		}
	}
	if last_o > 0 {
	tcc_define_symbol(s, c'__OPTIMIZE__', (voidptr(0)))
	}
	if linker_arg.size {
		r = linker_arg.data
		goto arg_err // id: 0x7fffc1f89688
	}
	*pargc = argc - arg_start
	*pargv = argv + arg_start
	if tool {
	return tool
	}
	if optind != noaction {
	return 0
	}
	if s.verbose == 2 {
	return 4
	}
	if s.verbose {
	return 3
	}
	return 1
}

fn tcc_set_options(s &TCCState, r &i8)  {
	argv := (voidptr(0))
	argc := 0
	args_parser_make_argv(r, &argc, &argv)
	tcc_parse_args(s, &argc, &argv, 0)
	dynarray_reset(&argv, &argc)
}

fn tcc_print_stats(s &TCCState, total_time u32)  {
	if total_time < 1 {
	total_time = 1
	}
	if total_bytes < 1 {
	total_bytes = 1
	}
	C.fprintf(C.stderr, c'* %d idents, %d lines, %d bytes\n* %0.3f s, %u lines/s, %0.1f MB/s\n', tok_ident - 256, total_lines, total_bytes, f64(total_time) / 1000, u32(total_lines) * 1000 / total_time, f64(total_bytes) / 1000 / total_time)
}

struct ArHdr { 
	ar_name [16]i8
	ar_date [12]i8
	ar_uid [6]i8
	ar_gid [6]i8
	ar_mode [8]i8
	ar_size [10]i8
	ar_fmag [2]i8
}
fn tcc_tool_ar(s1 &TCCState, argc int, argv &&u8) int {
	arhdr := ArHdr {
	ar_name: c'/               ', 
ar_date: c'            ', 
ar_uid: c'0     ', 
ar_gid: c'0     ', 
ar_mode: c'0       ', 
ar_size: c'          ', 
ar_fmag: c'`\n'
}
	
	arhdro := ArHdr {
	ar_name: c'                ', 
ar_date: c'            ', 
ar_uid: c'0     ', 
ar_gid: c'0     ', 
ar_mode: c'0       ', 
ar_size: c'          ', 
ar_fmag: c'`\n'
}
	
	fi := &C.FILE(0)
	fh := (voidptr(0))
fo := (voidptr(0))

	ehdr := &Elf64_Ehdr(0)
	shdr := &Elf64_Shdr(0)
	sym := &Elf64_Sym(0)
	i := 0
	fsize := 0
	i_lib := 0
	i_obj := 0
	
	buf := &i8(0)
	shstr := &i8(0)
	symtab := (voidptr(0))
strtab := (voidptr(0))

	symtabsize := 0
	anames := (voidptr(0))
	afpos := (voidptr(0))
	istrlen := 0
	strpos := 0
fpos := 0
funccnt := 0
funcmax := 0
	hofs := 0
	
	tfile := [260]i8{}
	stmp := [20]i8{}
	
	file := &i8(0)
	name := &i8(0)
	
	ret := 2
	ops_conflict := c'habdioptxN'
	verbose := 0
	i_lib = 0
	i_obj = 0
	for i = 1 ; i < argc ; i ++ {
		a := argv [i] 
		if *a == `-` && strstr(a, c'.') {
		ret = 1
		}
		if (*a == `-`) || (i == 1 && !strstr(a, c'.')) {
			if contains_any(a, ops_conflict) {
			ret = 1
			}
			if strstr(a, c'v') {
			verbose = 1
			}
		}
		else {
			if !i_lib {
			i_lib = i
			}
			else if !i_obj {
			i_obj = i
			}
		}
	}
	if !i_obj {
	ret = 1
	}
	if ret == 1 {
	return ar_usage(ret)
	}
	if (fh = C.fopen(argv [i_lib] , c'wb')) == (voidptr(0)) {
		C.fprintf(C.stderr, c"tcc: ar: can't open file %s \n", argv [i_lib] )
		goto the_end // id: 0x7fffc1f96f70
	}
	sprintf(tfile, c'%s.tmp', argv [i_lib] )
	if (fo = C.fopen(tfile, c'wb+')) == (voidptr(0)) {
		C.fprintf(C.stderr, c"tcc: ar: can't create temporary file %s\n", tfile)
		goto the_end // id: 0x7fffc1f96f70
	}
	funcmax = 250
	afpos = tcc_realloc((voidptr(0)), funcmax * sizeof*afpos)
	C.memcpy(&arhdro.ar_mode, c'100666', 6)
	for i_obj < argc {
		if *argv [i_obj]  == `-` {
			i_obj ++
			continue
			
		}
		if (fi = C.fopen(argv [i_obj] , c'rb')) == (voidptr(0)) {
			C.fprintf(C.stderr, c"tcc: ar: can't open file %s \n", argv [i_obj] )
			goto the_end // id: 0x7fffc1f96f70
		}
		if verbose {
		C.printf(c'a - %s\n', argv [i_obj] )
		}
		C.fseek(fi, 0, 2)
		fsize = C.ftell(fi)
		C.fseek(fi, 0, 0)
		buf = tcc_malloc(fsize + 1)
		C.fread(buf, fsize, 1, fi)
		C.fclose(fi)
		ehdr = &Elf64_Ehdr(buf)
		if ehdr.e_ident [4]  != 2 {
			C.fprintf(C.stderr, c'tcc: ar: Unsupported Elf Class: %s\n', argv [i_obj] )
			goto the_end // id: 0x7fffc1f96f70
		}
		shdr = &Elf64_Shdr((buf + ehdr.e_shoff + ehdr.e_shstrndx * ehdr.e_shentsize))
		shstr = &i8((buf + shdr.sh_offset))
		for i = 0 ; i < ehdr.e_shnum ; i ++ {
			shdr = &Elf64_Shdr((buf + ehdr.e_shoff + i * ehdr.e_shentsize))
			if !shdr.sh_offset {
			continue
			
			}
			if shdr.sh_type == 2 {
				symtab = &i8((buf + shdr.sh_offset))
				symtabsize = shdr.sh_size
			}
			if shdr.sh_type == 3 {
				if !C.strcmp(shstr + shdr.sh_name, c'.strtab') {
					strtab = &i8((buf + shdr.sh_offset))
				}
			}
		}
		if symtab && symtabsize {
			nsym := symtabsize / sizeof(Elf64_Sym)
			for i = 1 ; i < nsym ; i ++ {
				sym = &Elf64_Sym((symtab + i * sizeof(Elf64_Sym)))
				if sym.st_shndx && (sym.st_info == 16 || sym.st_info == 17 || sym.st_info == 18) {
					istrlen = C.strlen(strtab + sym.st_name) + 1
					anames = tcc_realloc(anames, strpos + istrlen)
					strcpy(anames + strpos, strtab + sym.st_name)
					strpos += istrlen
					if funccnt ++$ >= funcmax {
						funcmax += 250
						afpos = tcc_realloc(afpos, funcmax * sizeof*afpos)
					}
					afpos [funccnt]  = fpos
				}
			}
		}
		file = argv [i_obj] 
		for name = C.strchr(file, 0) ; name > file && name [-1]  != `/` && name [-1]  != `\\` ; name -- {
		0
		}
		istrlen = C.strlen(name)
		if istrlen >= sizeof(arhdro.ar_name) {
		istrlen = sizeof(arhdro.ar_name) - 1
		}
		C.memset(arhdro.ar_name, ` `, sizeof(arhdro.ar_name))
		C.memcpy(arhdro.ar_name, name, istrlen)
		arhdro.ar_name [istrlen]  = `/`
		sprintf(stmp, c'%-10d', fsize)
		C.memcpy(&arhdro.ar_size, stmp, 10)
		C.fwrite(&arhdro, sizeof(arhdro), 1, fo)
		C.fwrite(buf, fsize, 1, fo)
		tcc_free(buf)
		i_obj ++
		fpos += (fsize + sizeof(arhdro))
	}
	hofs = 8 + sizeof(arhdr) + strpos + (funccnt + 1) * sizeof(int)
	fpos = 0
	if (hofs & 1) {
	hofs ++ , 1
	fpos = hofs ++
	}
	C.fwrite(c'!<arch>\n', 8, 1, fh)
	sprintf(stmp, c'%-10d', int((strpos + (funccnt + 1) * sizeof(int))))
	C.memcpy(&arhdr.ar_size, stmp, 10)
	C.fwrite(&arhdr, sizeof(arhdr), 1, fh)
	afpos [0]  = le2belong(funccnt)
	for i = 1 ; i <= funccnt ; i ++ {
	afpos [i]  = le2belong(afpos [i]  + hofs)
	}
	C.fwrite(afpos, (funccnt + 1) * sizeof(int), 1, fh)
	C.fwrite(anames, strpos, 1, fh)
	if fpos {
	C.fwrite(c'', 1, 1, fh)
	}
	C.fseek(fo, 0, 2)
	fsize = C.ftell(fo)
	C.fseek(fo, 0, 0)
	buf = tcc_malloc(fsize + 1)
	C.fread(buf, fsize, 1, fo)
	C.fwrite(buf, fsize, 1, fh)
	tcc_free(buf)
	ret = 0
	// RRRREG the_end id=0x7fffc1f96f70
	the_end: 
	if anames {
	tcc_free(anames)
	}
	if afpos {
	tcc_free(afpos)
	}
	if fh {
	C.fclose(fh)
	}
	if fo {
	C.fclose(fo) , C.remove(tfile)
	}
	return ret
}

fn tcc_tool_cross(s &TCCState, argv &&u8, target int)  {
	program := [4096]i8{}
	a0 := argv [0] 
	prefix := tcc_basename(a0) - a0
	C.snprintf(program, sizeof(program), c'%.*s%s-tcc', prefix, a0, if target == 64{ c'x86_64' } else {c'i386'})
	if C.strcmp(a0, program) {
	execvp(argv [0]  = program, argv)
	}
	tcc_error(c"could not run '%s'", program)
}

fn gen_makedeps(s &TCCState, target &i8, filename &i8)  {
	depout := &C.FILE(0)
	buf := [1024]i8{}
	i := 0
	if !filename {
		C.snprintf(buf, sizeof(buf), c'%.*s.d', int((tcc_fileextension(target) - target)), target)
		filename = buf
	}
	if s.verbose {
	C.printf(c'<- %s\n', filename)
	}
	depout = C.fopen(filename, c'w')
	if !depout {
	tcc_error(c"could not open '%s'", filename)
	}
	C.fprintf(depout, c'%s: \\\n', target)
	for i = 0 ; i < s.nb_target_deps ; i ++ {
	C.fprintf(depout, c' %s \\\n', s.target_deps [i] )
	}
	C.fprintf(depout, c'\n')
	C.fclose(depout)
}

[export:'help']
const (
help   = c"Tiny C Compiler 0.9.27 - Copyright (C) 2001-2006 Fabrice Bellard\nUsage: tcc [options...] [-o outfile] [-c] infile(s)...\n       tcc [options...] -run infile [arguments...]\nGeneral options:\n  -c          compile only - generate an object file\n  -o outfile  set output filename\n  -run        run compiled source\n  -fflag      set or reset (with 'no-' prefix) 'flag' (see tcc -hh)\n  -std=c99    Conform to the ISO 1999 C standard (default).\n  -std=c11    Conform to the ISO 2011 C standard.\n  -Wwarning   set or reset (with 'no-' prefix) 'warning' (see tcc -hh)\n  -w          disable all warnings\n  -v -vv      show version, show search paths or loaded files\n  -h -hh      show this, show more help\n  -bench      show compilation statistics\n  -           use stdin pipe as infile\n  @listfile   read arguments from listfile\nPreprocessor options:\n  -Idir       add include path 'dir'\n  -Dsym[=val] define 'sym' with value 'val'\n  -Usym       undefine 'sym'\n  -E          preprocess only\nLinker options:\n  -Ldir       add library path 'dir'\n  -llib       link with dynamic or static library 'lib'\n  -r          generate (relocatable) object file\n  -shared     generate a shared library/dll\n  -rdynamic   export all global symbols to dynamic linker\n  -soname     set name for shared library to be used at runtime\n  -Wl,-opt[=val]  set linker option (see tcc -hh)\nDebugger options:\n  -g          generate runtime debug info\n  -b          compile with built-in memory and bounds checker (implies -g)\n  -bt N       show N callers in stack traces\nMisc. options:\n  -x[c|a|b|n] specify type of the next infile (C,ASM,BIN,NONE)\n  -nostdinc   do not use standard system include paths\n  -nostdlib   do not link with standard crt and libraries\n  -Bdir       set tcc's private include/library dir\n  -MD         generate dependency file for make\n  -MF file    specify dependency file name\n  -m32/64     defer to i386/x86_64 cross compiler\nTools:\n  create library  : tcc -ar [rcsv] lib.a files\n"
)

[export:'help2']
const (
help2   = c"Tiny C Compiler 0.9.27 - More Options\nSpecial options:\n  -P -P1                        with -E: no/alternative #line output\n  -dD -dM                       with -E: output #define directives\n  -pthread                      same as -D_REENTRANT and -lpthread\n  -On                           same as -D__OPTIMIZE__ for n > 0\n  -Wp,-opt                      same as -opt\n  -include file                 include 'file' above each input file\n  -isystem dir                  add 'dir' to system include path\n  -static                       link to static libraries (not recommended)\n  -dumpversion                  print version\n  -print-search-dirs            print search paths\n  -dt                           with -run/-E: auto-define 'test_...' macros\nIgnored options:\n  --param  -pedantic  -pipe  -s  -traditional\n-W... warnings:\n  all                           turn on some (*) warnings\n  error                         stop after first warning\n  unsupported                   warn about ignored options, pragmas, etc.\n  write-strings                 strings are const\n  implicit-function-declaration warn for missing prototype (*)\n-f[no-]... flags:\n  unsigned-char                 default char is unsigned\n  signed-char                   default char is signed\n  common                        use common section instead of bss\n  leading-underscore            decorate extern symbols\n  ms-extensions                 allow anonymous struct in struct\n  dollars-in-identifiers        allow '$' in C symbols\n-m... target specific options:\n  ms-bitfields                  use MSVC bitfield layout\n  no-sse                        disable floats on x86_64\n-Wl,... linker options:\n  -nostdlib                     do not link with standard crt/libs\n  -[no-]whole-archive           load lib(s) fully/only as needed\n  -export-all-symbols           same as -rdynamic\n  -export-dynamic               same as -rdynamic\n  -image-base= -Ttext=          set base address of executable\n  -section-alignment=           set section alignment in executable\n  -rpath=                       set dynamic library search path\n  -enable-new-dtags             set DT_RUNPATH instead of DT_RPATH\n  -soname=                      set DT_SONAME elf tag\n  -Bsymbolic                    set DT_SYMBOLIC elf tag\n  -oformat=[elf32/64-* binary]  set executable output format\n  -init= -fini= -as-needed -O   (ignored)\nPredefined macros:\n  tcc -E -dM - < /dev/null\nSee also the manual for more details.\n"
)

[export:'version']
const (
version   = c'tcc version 0.9.27 (x86_64 Linux)\n'
)

fn print_dirs(msg &i8, paths &&u8, nb_paths int)  {
	i := 0
	C.printf(c'%s:\n%s', msg, if nb_paths{ c'' } else {c'  -\n'})
	for i = 0 ; i < nb_paths ; i ++ {
	C.printf(c'  %s\n', paths [i] )
	}
}

fn print_search_dirs(s &TCCState)  {
	C.printf(c'install: %s\n', s.tcc_lib_path)
	print_dirs(c'include', s.sysinclude_paths, s.nb_sysinclude_paths)
	print_dirs(c'libraries', s.library_paths, s.nb_library_paths)
	C.printf(c'libtcc1:\n  %s/libtcc1.a\n', s.tcc_lib_path)
	print_dirs(c'crt', s.crt_paths, s.nb_crt_paths)
	C.printf(c'elfinterp:\n  %s\n', c'/lib64/ld-linux-x86-64.so.2')
}

fn set_environment(s &TCCState)  {
	path := &i8(0)
	path = getenv(c'C_INCLUDE_PATH')
	if path != (voidptr(0)) {
		tcc_add_sysinclude_path(s, path)
	}
	path = getenv(c'CPATH')
	if path != (voidptr(0)) {
		tcc_add_include_path(s, path)
	}
	path = getenv(c'LIBRARY_PATH')
	if path != (voidptr(0)) {
		tcc_add_library_path(s, path)
	}
}

fn default_outputfile(s &TCCState, first_file &i8) &i8 {
	buf := [1024]i8{}
	ext := &i8(0)
	name := c'a'
	if first_file && C.strcmp(first_file, c'-') {
	name = tcc_basename(first_file)
	}
	C.snprintf(buf, sizeof(buf), c'%s', name)
	ext = tcc_fileextension(buf)
	if s.output_type == 4 && !s.option_r && *ext {
	strcpy(ext, c'.o')
	}
	else { // 3
	strcpy(buf, c'a.out')
}
	return tcc_strdup(buf)
}

fn getclock_ms() u32 {
	tv := Timeval{}
	gettimeofday(&tv, (voidptr(0)))
	return tv.tv_sec * 1000 + (tv.tv_usec + 500) / 1000
}

fn main()  {
	s := &TCCState(0)
	ret := 0
	opt := 0
	n := 0
t := 0

	start_time := 0
	first_file := &i8(0)
	argc := 0
	argv := &&u8(0)
	ppfp := C.stdout
	// RRRREG redo id=0x7fffc1fabc30
	redo: 
	argc = argc0 , argv0
	argv = argc = argc0
	s = tcc_new()
	opt = tcc_parse_args(s, &argc, &argv, 1)
	if (n | t) == 0 {
		if opt == 1 {
		return 
		}
		if opt == 2 {
		return 
		}
		if opt == 32 || opt == 64 {
		tcc_tool_cross(s, argv, opt)
		}
		if s.verbose {
		C.printf(version)
		}
		if opt == 5 {
		return 
		}
		if opt == 3 {
		return 
		}
		if opt == 4 {
			set_environment(s)
			tcc_set_output_type(s, 1)
			print_search_dirs(s)
			return 
		}
		n = s.nb_files
		if n == 0 {
		tcc_error(c'no input files\n')
		}
		if s.output_type == 5 {
			if s.outfile && 0 != C.strcmp(c'-', s.outfile) {
				ppfp = C.fopen(s.outfile, c'w')
				if !ppfp {
				tcc_error(c"could not write '%s'", s.outfile)
				}
			}
		}
		else if s.output_type == 4 && !s.option_r {
			if s.nb_libraries {
			tcc_error(c'cannot specify libraries with -c')
			}
			if n > 1 && s.outfile {
			tcc_error(c'cannot specify output file with -c many files')
			}
		}
		else {
			if s.option_pthread {
				tcc_set_options(s, c'-lpthread')
				n = s.nb_files
			}
		}
		if s.do_bench {
		start_time = getclock_ms()
		}
	}
	set_environment(s)
	if s.output_type == 0 {
	s.output_type = 2
	}
	tcc_set_output_type(s, s.output_type)
	s.ppfp = ppfp
	if (s.output_type == 1 || s.output_type == 5) && (s.dflag & 16) {
	s.dflag |= if t{ 32 } else {0} , t ++$
	s.run_test = s.dflag |= if t{ 32 } else {0} , s.nb_files
	n = s.dflag |= if t{ 32 } else {0} , t ++$
	s.run_test = s.dflag |= if t{ 32 } else {0}
	}
	for first_file = (voidptr(0)) , 0
	ret = first_file = (voidptr(0)) ;  ;  {
		f := s.files [s.nb_files - n] 
		s.filetype = f.type_
		if f.type_ & 8 {
			if tcc_add_library_err(s, f.name) < 0 {
			ret = 1
			}
		}
		else {
			if 1 == s.verbose {
			C.printf(c'-> %s\n', f.name)
			}
			if !first_file {
			first_file = f.name
			}
			if tcc_add_file(s, f.name) < 0 {
			ret = 1
			}
		}
		if n --$ == 0 || ret || (s.output_type == 4 && !s.option_r) {
		break
		
		}
	}
	if s.run_test {
		t = 0
	}
	else if s.output_type == 5 {
		0
	}
	else if 0 == ret {
		if s.output_type == 1 {
			ret = tcc_run(s, argc, argv)
		}
		else {
			if !s.outfile {
			s.outfile = default_outputfile(s, first_file)
			}
			if tcc_output_file(s, s.outfile) {
			ret = 1
			}
			else if s.gen_deps {
			gen_makedeps(s, s.outfile, s.deps_outfile)
			}
		}
	}
	if s.do_bench && (n | t | ret) == 0 {
	tcc_print_stats(s, getclock_ms() - start_time)
	}
	tcc_delete(s)
	if ret == 0 && n {
	goto redo // id: 0x7fffc1fabc30
	}
	if t {
	goto redo // id: 0x7fffc1fabc30
	}
	if ppfp && ppfp != C.stdout {
	C.fclose(ppfp)
	}
	return 
}

