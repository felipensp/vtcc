@[translated]
module main

@[hidden; markused]
__global __dso_handle = unsafe { nil }
