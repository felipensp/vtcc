@[translated]
module main

__global dso_handle = unsafe { nil }
__global __dso_handle = &dso_handle
